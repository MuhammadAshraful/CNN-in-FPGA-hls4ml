
`include "dump_file_agent.svh"
`include "csv_file_dump.svh"
`include "sample_agent.svh"
`include "loop_sample_agent.svh"
`include "sample_manager.svh"
`include "nodf_module_interface.svh"
`include "nodf_module_monitor.svh"
`include "df_fifo_interface.svh"
`include "df_fifo_monitor.svh"
`include "df_process_interface.svh"
`include "df_process_monitor.svh"
`include "seq_loop_interface.svh"
`include "seq_loop_monitor.svh"
`include "upc_loop_interface.svh"
`include "upc_loop_monitor.svh"
`timescale 1ns/1ps

// top module for dataflow related monitors
module dataflow_monitor(
input logic clock,
input logic reset,
input logic finish
);

    df_fifo_intf fifo_intf_1(clock,reset);
    assign fifo_intf_1.rd_en = AESL_inst_myproject.layer2_out_U.if_read & AESL_inst_myproject.layer2_out_U.if_empty_n;
    assign fifo_intf_1.wr_en = AESL_inst_myproject.layer2_out_U.if_write & AESL_inst_myproject.layer2_out_U.if_full_n;
    assign fifo_intf_1.fifo_rd_block = 0;
    assign fifo_intf_1.fifo_wr_block = 0;
    assign fifo_intf_1.finish = finish;
    csv_file_dump fifo_csv_dumper_1;
    csv_file_dump cstatus_csv_dumper_1;
    df_fifo_monitor fifo_monitor_1;
    df_fifo_intf fifo_intf_2(clock,reset);
    assign fifo_intf_2.rd_en = AESL_inst_myproject.layer2_out_1_U.if_read & AESL_inst_myproject.layer2_out_1_U.if_empty_n;
    assign fifo_intf_2.wr_en = AESL_inst_myproject.layer2_out_1_U.if_write & AESL_inst_myproject.layer2_out_1_U.if_full_n;
    assign fifo_intf_2.fifo_rd_block = 0;
    assign fifo_intf_2.fifo_wr_block = 0;
    assign fifo_intf_2.finish = finish;
    csv_file_dump fifo_csv_dumper_2;
    csv_file_dump cstatus_csv_dumper_2;
    df_fifo_monitor fifo_monitor_2;
    df_fifo_intf fifo_intf_3(clock,reset);
    assign fifo_intf_3.rd_en = AESL_inst_myproject.layer2_out_2_U.if_read & AESL_inst_myproject.layer2_out_2_U.if_empty_n;
    assign fifo_intf_3.wr_en = AESL_inst_myproject.layer2_out_2_U.if_write & AESL_inst_myproject.layer2_out_2_U.if_full_n;
    assign fifo_intf_3.fifo_rd_block = 0;
    assign fifo_intf_3.fifo_wr_block = 0;
    assign fifo_intf_3.finish = finish;
    csv_file_dump fifo_csv_dumper_3;
    csv_file_dump cstatus_csv_dumper_3;
    df_fifo_monitor fifo_monitor_3;
    df_fifo_intf fifo_intf_4(clock,reset);
    assign fifo_intf_4.rd_en = AESL_inst_myproject.layer2_out_3_U.if_read & AESL_inst_myproject.layer2_out_3_U.if_empty_n;
    assign fifo_intf_4.wr_en = AESL_inst_myproject.layer2_out_3_U.if_write & AESL_inst_myproject.layer2_out_3_U.if_full_n;
    assign fifo_intf_4.fifo_rd_block = 0;
    assign fifo_intf_4.fifo_wr_block = 0;
    assign fifo_intf_4.finish = finish;
    csv_file_dump fifo_csv_dumper_4;
    csv_file_dump cstatus_csv_dumper_4;
    df_fifo_monitor fifo_monitor_4;
    df_fifo_intf fifo_intf_5(clock,reset);
    assign fifo_intf_5.rd_en = AESL_inst_myproject.layer2_out_4_U.if_read & AESL_inst_myproject.layer2_out_4_U.if_empty_n;
    assign fifo_intf_5.wr_en = AESL_inst_myproject.layer2_out_4_U.if_write & AESL_inst_myproject.layer2_out_4_U.if_full_n;
    assign fifo_intf_5.fifo_rd_block = 0;
    assign fifo_intf_5.fifo_wr_block = 0;
    assign fifo_intf_5.finish = finish;
    csv_file_dump fifo_csv_dumper_5;
    csv_file_dump cstatus_csv_dumper_5;
    df_fifo_monitor fifo_monitor_5;
    df_fifo_intf fifo_intf_6(clock,reset);
    assign fifo_intf_6.rd_en = AESL_inst_myproject.layer2_out_5_U.if_read & AESL_inst_myproject.layer2_out_5_U.if_empty_n;
    assign fifo_intf_6.wr_en = AESL_inst_myproject.layer2_out_5_U.if_write & AESL_inst_myproject.layer2_out_5_U.if_full_n;
    assign fifo_intf_6.fifo_rd_block = 0;
    assign fifo_intf_6.fifo_wr_block = 0;
    assign fifo_intf_6.finish = finish;
    csv_file_dump fifo_csv_dumper_6;
    csv_file_dump cstatus_csv_dumper_6;
    df_fifo_monitor fifo_monitor_6;
    df_fifo_intf fifo_intf_7(clock,reset);
    assign fifo_intf_7.rd_en = AESL_inst_myproject.layer2_out_6_U.if_read & AESL_inst_myproject.layer2_out_6_U.if_empty_n;
    assign fifo_intf_7.wr_en = AESL_inst_myproject.layer2_out_6_U.if_write & AESL_inst_myproject.layer2_out_6_U.if_full_n;
    assign fifo_intf_7.fifo_rd_block = 0;
    assign fifo_intf_7.fifo_wr_block = 0;
    assign fifo_intf_7.finish = finish;
    csv_file_dump fifo_csv_dumper_7;
    csv_file_dump cstatus_csv_dumper_7;
    df_fifo_monitor fifo_monitor_7;
    df_fifo_intf fifo_intf_8(clock,reset);
    assign fifo_intf_8.rd_en = AESL_inst_myproject.layer2_out_7_U.if_read & AESL_inst_myproject.layer2_out_7_U.if_empty_n;
    assign fifo_intf_8.wr_en = AESL_inst_myproject.layer2_out_7_U.if_write & AESL_inst_myproject.layer2_out_7_U.if_full_n;
    assign fifo_intf_8.fifo_rd_block = 0;
    assign fifo_intf_8.fifo_wr_block = 0;
    assign fifo_intf_8.finish = finish;
    csv_file_dump fifo_csv_dumper_8;
    csv_file_dump cstatus_csv_dumper_8;
    df_fifo_monitor fifo_monitor_8;
    df_fifo_intf fifo_intf_9(clock,reset);
    assign fifo_intf_9.rd_en = AESL_inst_myproject.layer2_out_8_U.if_read & AESL_inst_myproject.layer2_out_8_U.if_empty_n;
    assign fifo_intf_9.wr_en = AESL_inst_myproject.layer2_out_8_U.if_write & AESL_inst_myproject.layer2_out_8_U.if_full_n;
    assign fifo_intf_9.fifo_rd_block = 0;
    assign fifo_intf_9.fifo_wr_block = 0;
    assign fifo_intf_9.finish = finish;
    csv_file_dump fifo_csv_dumper_9;
    csv_file_dump cstatus_csv_dumper_9;
    df_fifo_monitor fifo_monitor_9;
    df_fifo_intf fifo_intf_10(clock,reset);
    assign fifo_intf_10.rd_en = AESL_inst_myproject.layer2_out_9_U.if_read & AESL_inst_myproject.layer2_out_9_U.if_empty_n;
    assign fifo_intf_10.wr_en = AESL_inst_myproject.layer2_out_9_U.if_write & AESL_inst_myproject.layer2_out_9_U.if_full_n;
    assign fifo_intf_10.fifo_rd_block = 0;
    assign fifo_intf_10.fifo_wr_block = 0;
    assign fifo_intf_10.finish = finish;
    csv_file_dump fifo_csv_dumper_10;
    csv_file_dump cstatus_csv_dumper_10;
    df_fifo_monitor fifo_monitor_10;
    df_fifo_intf fifo_intf_11(clock,reset);
    assign fifo_intf_11.rd_en = AESL_inst_myproject.layer2_out_10_U.if_read & AESL_inst_myproject.layer2_out_10_U.if_empty_n;
    assign fifo_intf_11.wr_en = AESL_inst_myproject.layer2_out_10_U.if_write & AESL_inst_myproject.layer2_out_10_U.if_full_n;
    assign fifo_intf_11.fifo_rd_block = 0;
    assign fifo_intf_11.fifo_wr_block = 0;
    assign fifo_intf_11.finish = finish;
    csv_file_dump fifo_csv_dumper_11;
    csv_file_dump cstatus_csv_dumper_11;
    df_fifo_monitor fifo_monitor_11;
    df_fifo_intf fifo_intf_12(clock,reset);
    assign fifo_intf_12.rd_en = AESL_inst_myproject.layer2_out_11_U.if_read & AESL_inst_myproject.layer2_out_11_U.if_empty_n;
    assign fifo_intf_12.wr_en = AESL_inst_myproject.layer2_out_11_U.if_write & AESL_inst_myproject.layer2_out_11_U.if_full_n;
    assign fifo_intf_12.fifo_rd_block = 0;
    assign fifo_intf_12.fifo_wr_block = 0;
    assign fifo_intf_12.finish = finish;
    csv_file_dump fifo_csv_dumper_12;
    csv_file_dump cstatus_csv_dumper_12;
    df_fifo_monitor fifo_monitor_12;
    df_fifo_intf fifo_intf_13(clock,reset);
    assign fifo_intf_13.rd_en = AESL_inst_myproject.layer2_out_12_U.if_read & AESL_inst_myproject.layer2_out_12_U.if_empty_n;
    assign fifo_intf_13.wr_en = AESL_inst_myproject.layer2_out_12_U.if_write & AESL_inst_myproject.layer2_out_12_U.if_full_n;
    assign fifo_intf_13.fifo_rd_block = 0;
    assign fifo_intf_13.fifo_wr_block = 0;
    assign fifo_intf_13.finish = finish;
    csv_file_dump fifo_csv_dumper_13;
    csv_file_dump cstatus_csv_dumper_13;
    df_fifo_monitor fifo_monitor_13;
    df_fifo_intf fifo_intf_14(clock,reset);
    assign fifo_intf_14.rd_en = AESL_inst_myproject.layer2_out_13_U.if_read & AESL_inst_myproject.layer2_out_13_U.if_empty_n;
    assign fifo_intf_14.wr_en = AESL_inst_myproject.layer2_out_13_U.if_write & AESL_inst_myproject.layer2_out_13_U.if_full_n;
    assign fifo_intf_14.fifo_rd_block = 0;
    assign fifo_intf_14.fifo_wr_block = 0;
    assign fifo_intf_14.finish = finish;
    csv_file_dump fifo_csv_dumper_14;
    csv_file_dump cstatus_csv_dumper_14;
    df_fifo_monitor fifo_monitor_14;
    df_fifo_intf fifo_intf_15(clock,reset);
    assign fifo_intf_15.rd_en = AESL_inst_myproject.layer2_out_14_U.if_read & AESL_inst_myproject.layer2_out_14_U.if_empty_n;
    assign fifo_intf_15.wr_en = AESL_inst_myproject.layer2_out_14_U.if_write & AESL_inst_myproject.layer2_out_14_U.if_full_n;
    assign fifo_intf_15.fifo_rd_block = 0;
    assign fifo_intf_15.fifo_wr_block = 0;
    assign fifo_intf_15.finish = finish;
    csv_file_dump fifo_csv_dumper_15;
    csv_file_dump cstatus_csv_dumper_15;
    df_fifo_monitor fifo_monitor_15;
    df_fifo_intf fifo_intf_16(clock,reset);
    assign fifo_intf_16.rd_en = AESL_inst_myproject.layer2_out_15_U.if_read & AESL_inst_myproject.layer2_out_15_U.if_empty_n;
    assign fifo_intf_16.wr_en = AESL_inst_myproject.layer2_out_15_U.if_write & AESL_inst_myproject.layer2_out_15_U.if_full_n;
    assign fifo_intf_16.fifo_rd_block = 0;
    assign fifo_intf_16.fifo_wr_block = 0;
    assign fifo_intf_16.finish = finish;
    csv_file_dump fifo_csv_dumper_16;
    csv_file_dump cstatus_csv_dumper_16;
    df_fifo_monitor fifo_monitor_16;
    df_fifo_intf fifo_intf_17(clock,reset);
    assign fifo_intf_17.rd_en = AESL_inst_myproject.layer2_out_16_U.if_read & AESL_inst_myproject.layer2_out_16_U.if_empty_n;
    assign fifo_intf_17.wr_en = AESL_inst_myproject.layer2_out_16_U.if_write & AESL_inst_myproject.layer2_out_16_U.if_full_n;
    assign fifo_intf_17.fifo_rd_block = 0;
    assign fifo_intf_17.fifo_wr_block = 0;
    assign fifo_intf_17.finish = finish;
    csv_file_dump fifo_csv_dumper_17;
    csv_file_dump cstatus_csv_dumper_17;
    df_fifo_monitor fifo_monitor_17;
    df_fifo_intf fifo_intf_18(clock,reset);
    assign fifo_intf_18.rd_en = AESL_inst_myproject.layer2_out_17_U.if_read & AESL_inst_myproject.layer2_out_17_U.if_empty_n;
    assign fifo_intf_18.wr_en = AESL_inst_myproject.layer2_out_17_U.if_write & AESL_inst_myproject.layer2_out_17_U.if_full_n;
    assign fifo_intf_18.fifo_rd_block = 0;
    assign fifo_intf_18.fifo_wr_block = 0;
    assign fifo_intf_18.finish = finish;
    csv_file_dump fifo_csv_dumper_18;
    csv_file_dump cstatus_csv_dumper_18;
    df_fifo_monitor fifo_monitor_18;
    df_fifo_intf fifo_intf_19(clock,reset);
    assign fifo_intf_19.rd_en = AESL_inst_myproject.layer2_out_18_U.if_read & AESL_inst_myproject.layer2_out_18_U.if_empty_n;
    assign fifo_intf_19.wr_en = AESL_inst_myproject.layer2_out_18_U.if_write & AESL_inst_myproject.layer2_out_18_U.if_full_n;
    assign fifo_intf_19.fifo_rd_block = 0;
    assign fifo_intf_19.fifo_wr_block = 0;
    assign fifo_intf_19.finish = finish;
    csv_file_dump fifo_csv_dumper_19;
    csv_file_dump cstatus_csv_dumper_19;
    df_fifo_monitor fifo_monitor_19;
    df_fifo_intf fifo_intf_20(clock,reset);
    assign fifo_intf_20.rd_en = AESL_inst_myproject.layer2_out_19_U.if_read & AESL_inst_myproject.layer2_out_19_U.if_empty_n;
    assign fifo_intf_20.wr_en = AESL_inst_myproject.layer2_out_19_U.if_write & AESL_inst_myproject.layer2_out_19_U.if_full_n;
    assign fifo_intf_20.fifo_rd_block = 0;
    assign fifo_intf_20.fifo_wr_block = 0;
    assign fifo_intf_20.finish = finish;
    csv_file_dump fifo_csv_dumper_20;
    csv_file_dump cstatus_csv_dumper_20;
    df_fifo_monitor fifo_monitor_20;
    df_fifo_intf fifo_intf_21(clock,reset);
    assign fifo_intf_21.rd_en = AESL_inst_myproject.layer2_out_20_U.if_read & AESL_inst_myproject.layer2_out_20_U.if_empty_n;
    assign fifo_intf_21.wr_en = AESL_inst_myproject.layer2_out_20_U.if_write & AESL_inst_myproject.layer2_out_20_U.if_full_n;
    assign fifo_intf_21.fifo_rd_block = 0;
    assign fifo_intf_21.fifo_wr_block = 0;
    assign fifo_intf_21.finish = finish;
    csv_file_dump fifo_csv_dumper_21;
    csv_file_dump cstatus_csv_dumper_21;
    df_fifo_monitor fifo_monitor_21;
    df_fifo_intf fifo_intf_22(clock,reset);
    assign fifo_intf_22.rd_en = AESL_inst_myproject.layer2_out_21_U.if_read & AESL_inst_myproject.layer2_out_21_U.if_empty_n;
    assign fifo_intf_22.wr_en = AESL_inst_myproject.layer2_out_21_U.if_write & AESL_inst_myproject.layer2_out_21_U.if_full_n;
    assign fifo_intf_22.fifo_rd_block = 0;
    assign fifo_intf_22.fifo_wr_block = 0;
    assign fifo_intf_22.finish = finish;
    csv_file_dump fifo_csv_dumper_22;
    csv_file_dump cstatus_csv_dumper_22;
    df_fifo_monitor fifo_monitor_22;
    df_fifo_intf fifo_intf_23(clock,reset);
    assign fifo_intf_23.rd_en = AESL_inst_myproject.layer2_out_22_U.if_read & AESL_inst_myproject.layer2_out_22_U.if_empty_n;
    assign fifo_intf_23.wr_en = AESL_inst_myproject.layer2_out_22_U.if_write & AESL_inst_myproject.layer2_out_22_U.if_full_n;
    assign fifo_intf_23.fifo_rd_block = 0;
    assign fifo_intf_23.fifo_wr_block = 0;
    assign fifo_intf_23.finish = finish;
    csv_file_dump fifo_csv_dumper_23;
    csv_file_dump cstatus_csv_dumper_23;
    df_fifo_monitor fifo_monitor_23;
    df_fifo_intf fifo_intf_24(clock,reset);
    assign fifo_intf_24.rd_en = AESL_inst_myproject.layer2_out_23_U.if_read & AESL_inst_myproject.layer2_out_23_U.if_empty_n;
    assign fifo_intf_24.wr_en = AESL_inst_myproject.layer2_out_23_U.if_write & AESL_inst_myproject.layer2_out_23_U.if_full_n;
    assign fifo_intf_24.fifo_rd_block = 0;
    assign fifo_intf_24.fifo_wr_block = 0;
    assign fifo_intf_24.finish = finish;
    csv_file_dump fifo_csv_dumper_24;
    csv_file_dump cstatus_csv_dumper_24;
    df_fifo_monitor fifo_monitor_24;
    df_fifo_intf fifo_intf_25(clock,reset);
    assign fifo_intf_25.rd_en = AESL_inst_myproject.layer2_out_24_U.if_read & AESL_inst_myproject.layer2_out_24_U.if_empty_n;
    assign fifo_intf_25.wr_en = AESL_inst_myproject.layer2_out_24_U.if_write & AESL_inst_myproject.layer2_out_24_U.if_full_n;
    assign fifo_intf_25.fifo_rd_block = 0;
    assign fifo_intf_25.fifo_wr_block = 0;
    assign fifo_intf_25.finish = finish;
    csv_file_dump fifo_csv_dumper_25;
    csv_file_dump cstatus_csv_dumper_25;
    df_fifo_monitor fifo_monitor_25;
    df_fifo_intf fifo_intf_26(clock,reset);
    assign fifo_intf_26.rd_en = AESL_inst_myproject.layer2_out_25_U.if_read & AESL_inst_myproject.layer2_out_25_U.if_empty_n;
    assign fifo_intf_26.wr_en = AESL_inst_myproject.layer2_out_25_U.if_write & AESL_inst_myproject.layer2_out_25_U.if_full_n;
    assign fifo_intf_26.fifo_rd_block = 0;
    assign fifo_intf_26.fifo_wr_block = 0;
    assign fifo_intf_26.finish = finish;
    csv_file_dump fifo_csv_dumper_26;
    csv_file_dump cstatus_csv_dumper_26;
    df_fifo_monitor fifo_monitor_26;
    df_fifo_intf fifo_intf_27(clock,reset);
    assign fifo_intf_27.rd_en = AESL_inst_myproject.layer2_out_26_U.if_read & AESL_inst_myproject.layer2_out_26_U.if_empty_n;
    assign fifo_intf_27.wr_en = AESL_inst_myproject.layer2_out_26_U.if_write & AESL_inst_myproject.layer2_out_26_U.if_full_n;
    assign fifo_intf_27.fifo_rd_block = 0;
    assign fifo_intf_27.fifo_wr_block = 0;
    assign fifo_intf_27.finish = finish;
    csv_file_dump fifo_csv_dumper_27;
    csv_file_dump cstatus_csv_dumper_27;
    df_fifo_monitor fifo_monitor_27;
    df_fifo_intf fifo_intf_28(clock,reset);
    assign fifo_intf_28.rd_en = AESL_inst_myproject.layer2_out_27_U.if_read & AESL_inst_myproject.layer2_out_27_U.if_empty_n;
    assign fifo_intf_28.wr_en = AESL_inst_myproject.layer2_out_27_U.if_write & AESL_inst_myproject.layer2_out_27_U.if_full_n;
    assign fifo_intf_28.fifo_rd_block = 0;
    assign fifo_intf_28.fifo_wr_block = 0;
    assign fifo_intf_28.finish = finish;
    csv_file_dump fifo_csv_dumper_28;
    csv_file_dump cstatus_csv_dumper_28;
    df_fifo_monitor fifo_monitor_28;
    df_fifo_intf fifo_intf_29(clock,reset);
    assign fifo_intf_29.rd_en = AESL_inst_myproject.layer2_out_28_U.if_read & AESL_inst_myproject.layer2_out_28_U.if_empty_n;
    assign fifo_intf_29.wr_en = AESL_inst_myproject.layer2_out_28_U.if_write & AESL_inst_myproject.layer2_out_28_U.if_full_n;
    assign fifo_intf_29.fifo_rd_block = 0;
    assign fifo_intf_29.fifo_wr_block = 0;
    assign fifo_intf_29.finish = finish;
    csv_file_dump fifo_csv_dumper_29;
    csv_file_dump cstatus_csv_dumper_29;
    df_fifo_monitor fifo_monitor_29;
    df_fifo_intf fifo_intf_30(clock,reset);
    assign fifo_intf_30.rd_en = AESL_inst_myproject.layer2_out_29_U.if_read & AESL_inst_myproject.layer2_out_29_U.if_empty_n;
    assign fifo_intf_30.wr_en = AESL_inst_myproject.layer2_out_29_U.if_write & AESL_inst_myproject.layer2_out_29_U.if_full_n;
    assign fifo_intf_30.fifo_rd_block = 0;
    assign fifo_intf_30.fifo_wr_block = 0;
    assign fifo_intf_30.finish = finish;
    csv_file_dump fifo_csv_dumper_30;
    csv_file_dump cstatus_csv_dumper_30;
    df_fifo_monitor fifo_monitor_30;
    df_fifo_intf fifo_intf_31(clock,reset);
    assign fifo_intf_31.rd_en = AESL_inst_myproject.layer2_out_30_U.if_read & AESL_inst_myproject.layer2_out_30_U.if_empty_n;
    assign fifo_intf_31.wr_en = AESL_inst_myproject.layer2_out_30_U.if_write & AESL_inst_myproject.layer2_out_30_U.if_full_n;
    assign fifo_intf_31.fifo_rd_block = 0;
    assign fifo_intf_31.fifo_wr_block = 0;
    assign fifo_intf_31.finish = finish;
    csv_file_dump fifo_csv_dumper_31;
    csv_file_dump cstatus_csv_dumper_31;
    df_fifo_monitor fifo_monitor_31;
    df_fifo_intf fifo_intf_32(clock,reset);
    assign fifo_intf_32.rd_en = AESL_inst_myproject.layer2_out_31_U.if_read & AESL_inst_myproject.layer2_out_31_U.if_empty_n;
    assign fifo_intf_32.wr_en = AESL_inst_myproject.layer2_out_31_U.if_write & AESL_inst_myproject.layer2_out_31_U.if_full_n;
    assign fifo_intf_32.fifo_rd_block = 0;
    assign fifo_intf_32.fifo_wr_block = 0;
    assign fifo_intf_32.finish = finish;
    csv_file_dump fifo_csv_dumper_32;
    csv_file_dump cstatus_csv_dumper_32;
    df_fifo_monitor fifo_monitor_32;
    df_fifo_intf fifo_intf_33(clock,reset);
    assign fifo_intf_33.rd_en = AESL_inst_myproject.layer2_out_32_U.if_read & AESL_inst_myproject.layer2_out_32_U.if_empty_n;
    assign fifo_intf_33.wr_en = AESL_inst_myproject.layer2_out_32_U.if_write & AESL_inst_myproject.layer2_out_32_U.if_full_n;
    assign fifo_intf_33.fifo_rd_block = 0;
    assign fifo_intf_33.fifo_wr_block = 0;
    assign fifo_intf_33.finish = finish;
    csv_file_dump fifo_csv_dumper_33;
    csv_file_dump cstatus_csv_dumper_33;
    df_fifo_monitor fifo_monitor_33;
    df_fifo_intf fifo_intf_34(clock,reset);
    assign fifo_intf_34.rd_en = AESL_inst_myproject.layer2_out_33_U.if_read & AESL_inst_myproject.layer2_out_33_U.if_empty_n;
    assign fifo_intf_34.wr_en = AESL_inst_myproject.layer2_out_33_U.if_write & AESL_inst_myproject.layer2_out_33_U.if_full_n;
    assign fifo_intf_34.fifo_rd_block = 0;
    assign fifo_intf_34.fifo_wr_block = 0;
    assign fifo_intf_34.finish = finish;
    csv_file_dump fifo_csv_dumper_34;
    csv_file_dump cstatus_csv_dumper_34;
    df_fifo_monitor fifo_monitor_34;
    df_fifo_intf fifo_intf_35(clock,reset);
    assign fifo_intf_35.rd_en = AESL_inst_myproject.layer2_out_34_U.if_read & AESL_inst_myproject.layer2_out_34_U.if_empty_n;
    assign fifo_intf_35.wr_en = AESL_inst_myproject.layer2_out_34_U.if_write & AESL_inst_myproject.layer2_out_34_U.if_full_n;
    assign fifo_intf_35.fifo_rd_block = 0;
    assign fifo_intf_35.fifo_wr_block = 0;
    assign fifo_intf_35.finish = finish;
    csv_file_dump fifo_csv_dumper_35;
    csv_file_dump cstatus_csv_dumper_35;
    df_fifo_monitor fifo_monitor_35;
    df_fifo_intf fifo_intf_36(clock,reset);
    assign fifo_intf_36.rd_en = AESL_inst_myproject.layer2_out_35_U.if_read & AESL_inst_myproject.layer2_out_35_U.if_empty_n;
    assign fifo_intf_36.wr_en = AESL_inst_myproject.layer2_out_35_U.if_write & AESL_inst_myproject.layer2_out_35_U.if_full_n;
    assign fifo_intf_36.fifo_rd_block = 0;
    assign fifo_intf_36.fifo_wr_block = 0;
    assign fifo_intf_36.finish = finish;
    csv_file_dump fifo_csv_dumper_36;
    csv_file_dump cstatus_csv_dumper_36;
    df_fifo_monitor fifo_monitor_36;
    df_fifo_intf fifo_intf_37(clock,reset);
    assign fifo_intf_37.rd_en = AESL_inst_myproject.layer2_out_36_U.if_read & AESL_inst_myproject.layer2_out_36_U.if_empty_n;
    assign fifo_intf_37.wr_en = AESL_inst_myproject.layer2_out_36_U.if_write & AESL_inst_myproject.layer2_out_36_U.if_full_n;
    assign fifo_intf_37.fifo_rd_block = 0;
    assign fifo_intf_37.fifo_wr_block = 0;
    assign fifo_intf_37.finish = finish;
    csv_file_dump fifo_csv_dumper_37;
    csv_file_dump cstatus_csv_dumper_37;
    df_fifo_monitor fifo_monitor_37;
    df_fifo_intf fifo_intf_38(clock,reset);
    assign fifo_intf_38.rd_en = AESL_inst_myproject.layer2_out_37_U.if_read & AESL_inst_myproject.layer2_out_37_U.if_empty_n;
    assign fifo_intf_38.wr_en = AESL_inst_myproject.layer2_out_37_U.if_write & AESL_inst_myproject.layer2_out_37_U.if_full_n;
    assign fifo_intf_38.fifo_rd_block = 0;
    assign fifo_intf_38.fifo_wr_block = 0;
    assign fifo_intf_38.finish = finish;
    csv_file_dump fifo_csv_dumper_38;
    csv_file_dump cstatus_csv_dumper_38;
    df_fifo_monitor fifo_monitor_38;
    df_fifo_intf fifo_intf_39(clock,reset);
    assign fifo_intf_39.rd_en = AESL_inst_myproject.layer2_out_38_U.if_read & AESL_inst_myproject.layer2_out_38_U.if_empty_n;
    assign fifo_intf_39.wr_en = AESL_inst_myproject.layer2_out_38_U.if_write & AESL_inst_myproject.layer2_out_38_U.if_full_n;
    assign fifo_intf_39.fifo_rd_block = 0;
    assign fifo_intf_39.fifo_wr_block = 0;
    assign fifo_intf_39.finish = finish;
    csv_file_dump fifo_csv_dumper_39;
    csv_file_dump cstatus_csv_dumper_39;
    df_fifo_monitor fifo_monitor_39;
    df_fifo_intf fifo_intf_40(clock,reset);
    assign fifo_intf_40.rd_en = AESL_inst_myproject.layer2_out_39_U.if_read & AESL_inst_myproject.layer2_out_39_U.if_empty_n;
    assign fifo_intf_40.wr_en = AESL_inst_myproject.layer2_out_39_U.if_write & AESL_inst_myproject.layer2_out_39_U.if_full_n;
    assign fifo_intf_40.fifo_rd_block = 0;
    assign fifo_intf_40.fifo_wr_block = 0;
    assign fifo_intf_40.finish = finish;
    csv_file_dump fifo_csv_dumper_40;
    csv_file_dump cstatus_csv_dumper_40;
    df_fifo_monitor fifo_monitor_40;
    df_fifo_intf fifo_intf_41(clock,reset);
    assign fifo_intf_41.rd_en = AESL_inst_myproject.layer2_out_40_U.if_read & AESL_inst_myproject.layer2_out_40_U.if_empty_n;
    assign fifo_intf_41.wr_en = AESL_inst_myproject.layer2_out_40_U.if_write & AESL_inst_myproject.layer2_out_40_U.if_full_n;
    assign fifo_intf_41.fifo_rd_block = 0;
    assign fifo_intf_41.fifo_wr_block = 0;
    assign fifo_intf_41.finish = finish;
    csv_file_dump fifo_csv_dumper_41;
    csv_file_dump cstatus_csv_dumper_41;
    df_fifo_monitor fifo_monitor_41;
    df_fifo_intf fifo_intf_42(clock,reset);
    assign fifo_intf_42.rd_en = AESL_inst_myproject.layer2_out_41_U.if_read & AESL_inst_myproject.layer2_out_41_U.if_empty_n;
    assign fifo_intf_42.wr_en = AESL_inst_myproject.layer2_out_41_U.if_write & AESL_inst_myproject.layer2_out_41_U.if_full_n;
    assign fifo_intf_42.fifo_rd_block = 0;
    assign fifo_intf_42.fifo_wr_block = 0;
    assign fifo_intf_42.finish = finish;
    csv_file_dump fifo_csv_dumper_42;
    csv_file_dump cstatus_csv_dumper_42;
    df_fifo_monitor fifo_monitor_42;
    df_fifo_intf fifo_intf_43(clock,reset);
    assign fifo_intf_43.rd_en = AESL_inst_myproject.layer2_out_42_U.if_read & AESL_inst_myproject.layer2_out_42_U.if_empty_n;
    assign fifo_intf_43.wr_en = AESL_inst_myproject.layer2_out_42_U.if_write & AESL_inst_myproject.layer2_out_42_U.if_full_n;
    assign fifo_intf_43.fifo_rd_block = 0;
    assign fifo_intf_43.fifo_wr_block = 0;
    assign fifo_intf_43.finish = finish;
    csv_file_dump fifo_csv_dumper_43;
    csv_file_dump cstatus_csv_dumper_43;
    df_fifo_monitor fifo_monitor_43;
    df_fifo_intf fifo_intf_44(clock,reset);
    assign fifo_intf_44.rd_en = AESL_inst_myproject.layer2_out_43_U.if_read & AESL_inst_myproject.layer2_out_43_U.if_empty_n;
    assign fifo_intf_44.wr_en = AESL_inst_myproject.layer2_out_43_U.if_write & AESL_inst_myproject.layer2_out_43_U.if_full_n;
    assign fifo_intf_44.fifo_rd_block = 0;
    assign fifo_intf_44.fifo_wr_block = 0;
    assign fifo_intf_44.finish = finish;
    csv_file_dump fifo_csv_dumper_44;
    csv_file_dump cstatus_csv_dumper_44;
    df_fifo_monitor fifo_monitor_44;
    df_fifo_intf fifo_intf_45(clock,reset);
    assign fifo_intf_45.rd_en = AESL_inst_myproject.layer2_out_44_U.if_read & AESL_inst_myproject.layer2_out_44_U.if_empty_n;
    assign fifo_intf_45.wr_en = AESL_inst_myproject.layer2_out_44_U.if_write & AESL_inst_myproject.layer2_out_44_U.if_full_n;
    assign fifo_intf_45.fifo_rd_block = 0;
    assign fifo_intf_45.fifo_wr_block = 0;
    assign fifo_intf_45.finish = finish;
    csv_file_dump fifo_csv_dumper_45;
    csv_file_dump cstatus_csv_dumper_45;
    df_fifo_monitor fifo_monitor_45;
    df_fifo_intf fifo_intf_46(clock,reset);
    assign fifo_intf_46.rd_en = AESL_inst_myproject.layer2_out_45_U.if_read & AESL_inst_myproject.layer2_out_45_U.if_empty_n;
    assign fifo_intf_46.wr_en = AESL_inst_myproject.layer2_out_45_U.if_write & AESL_inst_myproject.layer2_out_45_U.if_full_n;
    assign fifo_intf_46.fifo_rd_block = 0;
    assign fifo_intf_46.fifo_wr_block = 0;
    assign fifo_intf_46.finish = finish;
    csv_file_dump fifo_csv_dumper_46;
    csv_file_dump cstatus_csv_dumper_46;
    df_fifo_monitor fifo_monitor_46;
    df_fifo_intf fifo_intf_47(clock,reset);
    assign fifo_intf_47.rd_en = AESL_inst_myproject.layer2_out_46_U.if_read & AESL_inst_myproject.layer2_out_46_U.if_empty_n;
    assign fifo_intf_47.wr_en = AESL_inst_myproject.layer2_out_46_U.if_write & AESL_inst_myproject.layer2_out_46_U.if_full_n;
    assign fifo_intf_47.fifo_rd_block = 0;
    assign fifo_intf_47.fifo_wr_block = 0;
    assign fifo_intf_47.finish = finish;
    csv_file_dump fifo_csv_dumper_47;
    csv_file_dump cstatus_csv_dumper_47;
    df_fifo_monitor fifo_monitor_47;
    df_fifo_intf fifo_intf_48(clock,reset);
    assign fifo_intf_48.rd_en = AESL_inst_myproject.layer2_out_47_U.if_read & AESL_inst_myproject.layer2_out_47_U.if_empty_n;
    assign fifo_intf_48.wr_en = AESL_inst_myproject.layer2_out_47_U.if_write & AESL_inst_myproject.layer2_out_47_U.if_full_n;
    assign fifo_intf_48.fifo_rd_block = 0;
    assign fifo_intf_48.fifo_wr_block = 0;
    assign fifo_intf_48.finish = finish;
    csv_file_dump fifo_csv_dumper_48;
    csv_file_dump cstatus_csv_dumper_48;
    df_fifo_monitor fifo_monitor_48;
    df_fifo_intf fifo_intf_49(clock,reset);
    assign fifo_intf_49.rd_en = AESL_inst_myproject.layer2_out_48_U.if_read & AESL_inst_myproject.layer2_out_48_U.if_empty_n;
    assign fifo_intf_49.wr_en = AESL_inst_myproject.layer2_out_48_U.if_write & AESL_inst_myproject.layer2_out_48_U.if_full_n;
    assign fifo_intf_49.fifo_rd_block = 0;
    assign fifo_intf_49.fifo_wr_block = 0;
    assign fifo_intf_49.finish = finish;
    csv_file_dump fifo_csv_dumper_49;
    csv_file_dump cstatus_csv_dumper_49;
    df_fifo_monitor fifo_monitor_49;
    df_fifo_intf fifo_intf_50(clock,reset);
    assign fifo_intf_50.rd_en = AESL_inst_myproject.layer2_out_49_U.if_read & AESL_inst_myproject.layer2_out_49_U.if_empty_n;
    assign fifo_intf_50.wr_en = AESL_inst_myproject.layer2_out_49_U.if_write & AESL_inst_myproject.layer2_out_49_U.if_full_n;
    assign fifo_intf_50.fifo_rd_block = 0;
    assign fifo_intf_50.fifo_wr_block = 0;
    assign fifo_intf_50.finish = finish;
    csv_file_dump fifo_csv_dumper_50;
    csv_file_dump cstatus_csv_dumper_50;
    df_fifo_monitor fifo_monitor_50;
    df_fifo_intf fifo_intf_51(clock,reset);
    assign fifo_intf_51.rd_en = AESL_inst_myproject.layer2_out_50_U.if_read & AESL_inst_myproject.layer2_out_50_U.if_empty_n;
    assign fifo_intf_51.wr_en = AESL_inst_myproject.layer2_out_50_U.if_write & AESL_inst_myproject.layer2_out_50_U.if_full_n;
    assign fifo_intf_51.fifo_rd_block = 0;
    assign fifo_intf_51.fifo_wr_block = 0;
    assign fifo_intf_51.finish = finish;
    csv_file_dump fifo_csv_dumper_51;
    csv_file_dump cstatus_csv_dumper_51;
    df_fifo_monitor fifo_monitor_51;
    df_fifo_intf fifo_intf_52(clock,reset);
    assign fifo_intf_52.rd_en = AESL_inst_myproject.layer2_out_51_U.if_read & AESL_inst_myproject.layer2_out_51_U.if_empty_n;
    assign fifo_intf_52.wr_en = AESL_inst_myproject.layer2_out_51_U.if_write & AESL_inst_myproject.layer2_out_51_U.if_full_n;
    assign fifo_intf_52.fifo_rd_block = 0;
    assign fifo_intf_52.fifo_wr_block = 0;
    assign fifo_intf_52.finish = finish;
    csv_file_dump fifo_csv_dumper_52;
    csv_file_dump cstatus_csv_dumper_52;
    df_fifo_monitor fifo_monitor_52;
    df_fifo_intf fifo_intf_53(clock,reset);
    assign fifo_intf_53.rd_en = AESL_inst_myproject.layer2_out_52_U.if_read & AESL_inst_myproject.layer2_out_52_U.if_empty_n;
    assign fifo_intf_53.wr_en = AESL_inst_myproject.layer2_out_52_U.if_write & AESL_inst_myproject.layer2_out_52_U.if_full_n;
    assign fifo_intf_53.fifo_rd_block = 0;
    assign fifo_intf_53.fifo_wr_block = 0;
    assign fifo_intf_53.finish = finish;
    csv_file_dump fifo_csv_dumper_53;
    csv_file_dump cstatus_csv_dumper_53;
    df_fifo_monitor fifo_monitor_53;
    df_fifo_intf fifo_intf_54(clock,reset);
    assign fifo_intf_54.rd_en = AESL_inst_myproject.layer2_out_53_U.if_read & AESL_inst_myproject.layer2_out_53_U.if_empty_n;
    assign fifo_intf_54.wr_en = AESL_inst_myproject.layer2_out_53_U.if_write & AESL_inst_myproject.layer2_out_53_U.if_full_n;
    assign fifo_intf_54.fifo_rd_block = 0;
    assign fifo_intf_54.fifo_wr_block = 0;
    assign fifo_intf_54.finish = finish;
    csv_file_dump fifo_csv_dumper_54;
    csv_file_dump cstatus_csv_dumper_54;
    df_fifo_monitor fifo_monitor_54;
    df_fifo_intf fifo_intf_55(clock,reset);
    assign fifo_intf_55.rd_en = AESL_inst_myproject.layer2_out_54_U.if_read & AESL_inst_myproject.layer2_out_54_U.if_empty_n;
    assign fifo_intf_55.wr_en = AESL_inst_myproject.layer2_out_54_U.if_write & AESL_inst_myproject.layer2_out_54_U.if_full_n;
    assign fifo_intf_55.fifo_rd_block = 0;
    assign fifo_intf_55.fifo_wr_block = 0;
    assign fifo_intf_55.finish = finish;
    csv_file_dump fifo_csv_dumper_55;
    csv_file_dump cstatus_csv_dumper_55;
    df_fifo_monitor fifo_monitor_55;
    df_fifo_intf fifo_intf_56(clock,reset);
    assign fifo_intf_56.rd_en = AESL_inst_myproject.layer2_out_55_U.if_read & AESL_inst_myproject.layer2_out_55_U.if_empty_n;
    assign fifo_intf_56.wr_en = AESL_inst_myproject.layer2_out_55_U.if_write & AESL_inst_myproject.layer2_out_55_U.if_full_n;
    assign fifo_intf_56.fifo_rd_block = 0;
    assign fifo_intf_56.fifo_wr_block = 0;
    assign fifo_intf_56.finish = finish;
    csv_file_dump fifo_csv_dumper_56;
    csv_file_dump cstatus_csv_dumper_56;
    df_fifo_monitor fifo_monitor_56;
    df_fifo_intf fifo_intf_57(clock,reset);
    assign fifo_intf_57.rd_en = AESL_inst_myproject.layer2_out_56_U.if_read & AESL_inst_myproject.layer2_out_56_U.if_empty_n;
    assign fifo_intf_57.wr_en = AESL_inst_myproject.layer2_out_56_U.if_write & AESL_inst_myproject.layer2_out_56_U.if_full_n;
    assign fifo_intf_57.fifo_rd_block = 0;
    assign fifo_intf_57.fifo_wr_block = 0;
    assign fifo_intf_57.finish = finish;
    csv_file_dump fifo_csv_dumper_57;
    csv_file_dump cstatus_csv_dumper_57;
    df_fifo_monitor fifo_monitor_57;
    df_fifo_intf fifo_intf_58(clock,reset);
    assign fifo_intf_58.rd_en = AESL_inst_myproject.layer2_out_57_U.if_read & AESL_inst_myproject.layer2_out_57_U.if_empty_n;
    assign fifo_intf_58.wr_en = AESL_inst_myproject.layer2_out_57_U.if_write & AESL_inst_myproject.layer2_out_57_U.if_full_n;
    assign fifo_intf_58.fifo_rd_block = 0;
    assign fifo_intf_58.fifo_wr_block = 0;
    assign fifo_intf_58.finish = finish;
    csv_file_dump fifo_csv_dumper_58;
    csv_file_dump cstatus_csv_dumper_58;
    df_fifo_monitor fifo_monitor_58;
    df_fifo_intf fifo_intf_59(clock,reset);
    assign fifo_intf_59.rd_en = AESL_inst_myproject.layer2_out_58_U.if_read & AESL_inst_myproject.layer2_out_58_U.if_empty_n;
    assign fifo_intf_59.wr_en = AESL_inst_myproject.layer2_out_58_U.if_write & AESL_inst_myproject.layer2_out_58_U.if_full_n;
    assign fifo_intf_59.fifo_rd_block = 0;
    assign fifo_intf_59.fifo_wr_block = 0;
    assign fifo_intf_59.finish = finish;
    csv_file_dump fifo_csv_dumper_59;
    csv_file_dump cstatus_csv_dumper_59;
    df_fifo_monitor fifo_monitor_59;
    df_fifo_intf fifo_intf_60(clock,reset);
    assign fifo_intf_60.rd_en = AESL_inst_myproject.layer2_out_59_U.if_read & AESL_inst_myproject.layer2_out_59_U.if_empty_n;
    assign fifo_intf_60.wr_en = AESL_inst_myproject.layer2_out_59_U.if_write & AESL_inst_myproject.layer2_out_59_U.if_full_n;
    assign fifo_intf_60.fifo_rd_block = 0;
    assign fifo_intf_60.fifo_wr_block = 0;
    assign fifo_intf_60.finish = finish;
    csv_file_dump fifo_csv_dumper_60;
    csv_file_dump cstatus_csv_dumper_60;
    df_fifo_monitor fifo_monitor_60;
    df_fifo_intf fifo_intf_61(clock,reset);
    assign fifo_intf_61.rd_en = AESL_inst_myproject.layer2_out_60_U.if_read & AESL_inst_myproject.layer2_out_60_U.if_empty_n;
    assign fifo_intf_61.wr_en = AESL_inst_myproject.layer2_out_60_U.if_write & AESL_inst_myproject.layer2_out_60_U.if_full_n;
    assign fifo_intf_61.fifo_rd_block = 0;
    assign fifo_intf_61.fifo_wr_block = 0;
    assign fifo_intf_61.finish = finish;
    csv_file_dump fifo_csv_dumper_61;
    csv_file_dump cstatus_csv_dumper_61;
    df_fifo_monitor fifo_monitor_61;
    df_fifo_intf fifo_intf_62(clock,reset);
    assign fifo_intf_62.rd_en = AESL_inst_myproject.layer2_out_61_U.if_read & AESL_inst_myproject.layer2_out_61_U.if_empty_n;
    assign fifo_intf_62.wr_en = AESL_inst_myproject.layer2_out_61_U.if_write & AESL_inst_myproject.layer2_out_61_U.if_full_n;
    assign fifo_intf_62.fifo_rd_block = 0;
    assign fifo_intf_62.fifo_wr_block = 0;
    assign fifo_intf_62.finish = finish;
    csv_file_dump fifo_csv_dumper_62;
    csv_file_dump cstatus_csv_dumper_62;
    df_fifo_monitor fifo_monitor_62;
    df_fifo_intf fifo_intf_63(clock,reset);
    assign fifo_intf_63.rd_en = AESL_inst_myproject.layer2_out_62_U.if_read & AESL_inst_myproject.layer2_out_62_U.if_empty_n;
    assign fifo_intf_63.wr_en = AESL_inst_myproject.layer2_out_62_U.if_write & AESL_inst_myproject.layer2_out_62_U.if_full_n;
    assign fifo_intf_63.fifo_rd_block = 0;
    assign fifo_intf_63.fifo_wr_block = 0;
    assign fifo_intf_63.finish = finish;
    csv_file_dump fifo_csv_dumper_63;
    csv_file_dump cstatus_csv_dumper_63;
    df_fifo_monitor fifo_monitor_63;
    df_fifo_intf fifo_intf_64(clock,reset);
    assign fifo_intf_64.rd_en = AESL_inst_myproject.layer2_out_63_U.if_read & AESL_inst_myproject.layer2_out_63_U.if_empty_n;
    assign fifo_intf_64.wr_en = AESL_inst_myproject.layer2_out_63_U.if_write & AESL_inst_myproject.layer2_out_63_U.if_full_n;
    assign fifo_intf_64.fifo_rd_block = 0;
    assign fifo_intf_64.fifo_wr_block = 0;
    assign fifo_intf_64.finish = finish;
    csv_file_dump fifo_csv_dumper_64;
    csv_file_dump cstatus_csv_dumper_64;
    df_fifo_monitor fifo_monitor_64;
    df_fifo_intf fifo_intf_65(clock,reset);
    assign fifo_intf_65.rd_en = AESL_inst_myproject.layer2_out_64_U.if_read & AESL_inst_myproject.layer2_out_64_U.if_empty_n;
    assign fifo_intf_65.wr_en = AESL_inst_myproject.layer2_out_64_U.if_write & AESL_inst_myproject.layer2_out_64_U.if_full_n;
    assign fifo_intf_65.fifo_rd_block = 0;
    assign fifo_intf_65.fifo_wr_block = 0;
    assign fifo_intf_65.finish = finish;
    csv_file_dump fifo_csv_dumper_65;
    csv_file_dump cstatus_csv_dumper_65;
    df_fifo_monitor fifo_monitor_65;
    df_fifo_intf fifo_intf_66(clock,reset);
    assign fifo_intf_66.rd_en = AESL_inst_myproject.layer2_out_65_U.if_read & AESL_inst_myproject.layer2_out_65_U.if_empty_n;
    assign fifo_intf_66.wr_en = AESL_inst_myproject.layer2_out_65_U.if_write & AESL_inst_myproject.layer2_out_65_U.if_full_n;
    assign fifo_intf_66.fifo_rd_block = 0;
    assign fifo_intf_66.fifo_wr_block = 0;
    assign fifo_intf_66.finish = finish;
    csv_file_dump fifo_csv_dumper_66;
    csv_file_dump cstatus_csv_dumper_66;
    df_fifo_monitor fifo_monitor_66;
    df_fifo_intf fifo_intf_67(clock,reset);
    assign fifo_intf_67.rd_en = AESL_inst_myproject.layer2_out_66_U.if_read & AESL_inst_myproject.layer2_out_66_U.if_empty_n;
    assign fifo_intf_67.wr_en = AESL_inst_myproject.layer2_out_66_U.if_write & AESL_inst_myproject.layer2_out_66_U.if_full_n;
    assign fifo_intf_67.fifo_rd_block = 0;
    assign fifo_intf_67.fifo_wr_block = 0;
    assign fifo_intf_67.finish = finish;
    csv_file_dump fifo_csv_dumper_67;
    csv_file_dump cstatus_csv_dumper_67;
    df_fifo_monitor fifo_monitor_67;
    df_fifo_intf fifo_intf_68(clock,reset);
    assign fifo_intf_68.rd_en = AESL_inst_myproject.layer2_out_67_U.if_read & AESL_inst_myproject.layer2_out_67_U.if_empty_n;
    assign fifo_intf_68.wr_en = AESL_inst_myproject.layer2_out_67_U.if_write & AESL_inst_myproject.layer2_out_67_U.if_full_n;
    assign fifo_intf_68.fifo_rd_block = 0;
    assign fifo_intf_68.fifo_wr_block = 0;
    assign fifo_intf_68.finish = finish;
    csv_file_dump fifo_csv_dumper_68;
    csv_file_dump cstatus_csv_dumper_68;
    df_fifo_monitor fifo_monitor_68;
    df_fifo_intf fifo_intf_69(clock,reset);
    assign fifo_intf_69.rd_en = AESL_inst_myproject.layer2_out_68_U.if_read & AESL_inst_myproject.layer2_out_68_U.if_empty_n;
    assign fifo_intf_69.wr_en = AESL_inst_myproject.layer2_out_68_U.if_write & AESL_inst_myproject.layer2_out_68_U.if_full_n;
    assign fifo_intf_69.fifo_rd_block = 0;
    assign fifo_intf_69.fifo_wr_block = 0;
    assign fifo_intf_69.finish = finish;
    csv_file_dump fifo_csv_dumper_69;
    csv_file_dump cstatus_csv_dumper_69;
    df_fifo_monitor fifo_monitor_69;
    df_fifo_intf fifo_intf_70(clock,reset);
    assign fifo_intf_70.rd_en = AESL_inst_myproject.layer2_out_69_U.if_read & AESL_inst_myproject.layer2_out_69_U.if_empty_n;
    assign fifo_intf_70.wr_en = AESL_inst_myproject.layer2_out_69_U.if_write & AESL_inst_myproject.layer2_out_69_U.if_full_n;
    assign fifo_intf_70.fifo_rd_block = 0;
    assign fifo_intf_70.fifo_wr_block = 0;
    assign fifo_intf_70.finish = finish;
    csv_file_dump fifo_csv_dumper_70;
    csv_file_dump cstatus_csv_dumper_70;
    df_fifo_monitor fifo_monitor_70;
    df_fifo_intf fifo_intf_71(clock,reset);
    assign fifo_intf_71.rd_en = AESL_inst_myproject.layer2_out_70_U.if_read & AESL_inst_myproject.layer2_out_70_U.if_empty_n;
    assign fifo_intf_71.wr_en = AESL_inst_myproject.layer2_out_70_U.if_write & AESL_inst_myproject.layer2_out_70_U.if_full_n;
    assign fifo_intf_71.fifo_rd_block = 0;
    assign fifo_intf_71.fifo_wr_block = 0;
    assign fifo_intf_71.finish = finish;
    csv_file_dump fifo_csv_dumper_71;
    csv_file_dump cstatus_csv_dumper_71;
    df_fifo_monitor fifo_monitor_71;
    df_fifo_intf fifo_intf_72(clock,reset);
    assign fifo_intf_72.rd_en = AESL_inst_myproject.layer2_out_71_U.if_read & AESL_inst_myproject.layer2_out_71_U.if_empty_n;
    assign fifo_intf_72.wr_en = AESL_inst_myproject.layer2_out_71_U.if_write & AESL_inst_myproject.layer2_out_71_U.if_full_n;
    assign fifo_intf_72.fifo_rd_block = 0;
    assign fifo_intf_72.fifo_wr_block = 0;
    assign fifo_intf_72.finish = finish;
    csv_file_dump fifo_csv_dumper_72;
    csv_file_dump cstatus_csv_dumper_72;
    df_fifo_monitor fifo_monitor_72;
    df_fifo_intf fifo_intf_73(clock,reset);
    assign fifo_intf_73.rd_en = AESL_inst_myproject.layer2_out_72_U.if_read & AESL_inst_myproject.layer2_out_72_U.if_empty_n;
    assign fifo_intf_73.wr_en = AESL_inst_myproject.layer2_out_72_U.if_write & AESL_inst_myproject.layer2_out_72_U.if_full_n;
    assign fifo_intf_73.fifo_rd_block = 0;
    assign fifo_intf_73.fifo_wr_block = 0;
    assign fifo_intf_73.finish = finish;
    csv_file_dump fifo_csv_dumper_73;
    csv_file_dump cstatus_csv_dumper_73;
    df_fifo_monitor fifo_monitor_73;
    df_fifo_intf fifo_intf_74(clock,reset);
    assign fifo_intf_74.rd_en = AESL_inst_myproject.layer2_out_73_U.if_read & AESL_inst_myproject.layer2_out_73_U.if_empty_n;
    assign fifo_intf_74.wr_en = AESL_inst_myproject.layer2_out_73_U.if_write & AESL_inst_myproject.layer2_out_73_U.if_full_n;
    assign fifo_intf_74.fifo_rd_block = 0;
    assign fifo_intf_74.fifo_wr_block = 0;
    assign fifo_intf_74.finish = finish;
    csv_file_dump fifo_csv_dumper_74;
    csv_file_dump cstatus_csv_dumper_74;
    df_fifo_monitor fifo_monitor_74;
    df_fifo_intf fifo_intf_75(clock,reset);
    assign fifo_intf_75.rd_en = AESL_inst_myproject.layer2_out_74_U.if_read & AESL_inst_myproject.layer2_out_74_U.if_empty_n;
    assign fifo_intf_75.wr_en = AESL_inst_myproject.layer2_out_74_U.if_write & AESL_inst_myproject.layer2_out_74_U.if_full_n;
    assign fifo_intf_75.fifo_rd_block = 0;
    assign fifo_intf_75.fifo_wr_block = 0;
    assign fifo_intf_75.finish = finish;
    csv_file_dump fifo_csv_dumper_75;
    csv_file_dump cstatus_csv_dumper_75;
    df_fifo_monitor fifo_monitor_75;
    df_fifo_intf fifo_intf_76(clock,reset);
    assign fifo_intf_76.rd_en = AESL_inst_myproject.layer2_out_75_U.if_read & AESL_inst_myproject.layer2_out_75_U.if_empty_n;
    assign fifo_intf_76.wr_en = AESL_inst_myproject.layer2_out_75_U.if_write & AESL_inst_myproject.layer2_out_75_U.if_full_n;
    assign fifo_intf_76.fifo_rd_block = 0;
    assign fifo_intf_76.fifo_wr_block = 0;
    assign fifo_intf_76.finish = finish;
    csv_file_dump fifo_csv_dumper_76;
    csv_file_dump cstatus_csv_dumper_76;
    df_fifo_monitor fifo_monitor_76;
    df_fifo_intf fifo_intf_77(clock,reset);
    assign fifo_intf_77.rd_en = AESL_inst_myproject.layer2_out_76_U.if_read & AESL_inst_myproject.layer2_out_76_U.if_empty_n;
    assign fifo_intf_77.wr_en = AESL_inst_myproject.layer2_out_76_U.if_write & AESL_inst_myproject.layer2_out_76_U.if_full_n;
    assign fifo_intf_77.fifo_rd_block = 0;
    assign fifo_intf_77.fifo_wr_block = 0;
    assign fifo_intf_77.finish = finish;
    csv_file_dump fifo_csv_dumper_77;
    csv_file_dump cstatus_csv_dumper_77;
    df_fifo_monitor fifo_monitor_77;
    df_fifo_intf fifo_intf_78(clock,reset);
    assign fifo_intf_78.rd_en = AESL_inst_myproject.layer2_out_77_U.if_read & AESL_inst_myproject.layer2_out_77_U.if_empty_n;
    assign fifo_intf_78.wr_en = AESL_inst_myproject.layer2_out_77_U.if_write & AESL_inst_myproject.layer2_out_77_U.if_full_n;
    assign fifo_intf_78.fifo_rd_block = 0;
    assign fifo_intf_78.fifo_wr_block = 0;
    assign fifo_intf_78.finish = finish;
    csv_file_dump fifo_csv_dumper_78;
    csv_file_dump cstatus_csv_dumper_78;
    df_fifo_monitor fifo_monitor_78;
    df_fifo_intf fifo_intf_79(clock,reset);
    assign fifo_intf_79.rd_en = AESL_inst_myproject.layer2_out_78_U.if_read & AESL_inst_myproject.layer2_out_78_U.if_empty_n;
    assign fifo_intf_79.wr_en = AESL_inst_myproject.layer2_out_78_U.if_write & AESL_inst_myproject.layer2_out_78_U.if_full_n;
    assign fifo_intf_79.fifo_rd_block = 0;
    assign fifo_intf_79.fifo_wr_block = 0;
    assign fifo_intf_79.finish = finish;
    csv_file_dump fifo_csv_dumper_79;
    csv_file_dump cstatus_csv_dumper_79;
    df_fifo_monitor fifo_monitor_79;
    df_fifo_intf fifo_intf_80(clock,reset);
    assign fifo_intf_80.rd_en = AESL_inst_myproject.layer2_out_79_U.if_read & AESL_inst_myproject.layer2_out_79_U.if_empty_n;
    assign fifo_intf_80.wr_en = AESL_inst_myproject.layer2_out_79_U.if_write & AESL_inst_myproject.layer2_out_79_U.if_full_n;
    assign fifo_intf_80.fifo_rd_block = 0;
    assign fifo_intf_80.fifo_wr_block = 0;
    assign fifo_intf_80.finish = finish;
    csv_file_dump fifo_csv_dumper_80;
    csv_file_dump cstatus_csv_dumper_80;
    df_fifo_monitor fifo_monitor_80;
    df_fifo_intf fifo_intf_81(clock,reset);
    assign fifo_intf_81.rd_en = AESL_inst_myproject.layer2_out_80_U.if_read & AESL_inst_myproject.layer2_out_80_U.if_empty_n;
    assign fifo_intf_81.wr_en = AESL_inst_myproject.layer2_out_80_U.if_write & AESL_inst_myproject.layer2_out_80_U.if_full_n;
    assign fifo_intf_81.fifo_rd_block = 0;
    assign fifo_intf_81.fifo_wr_block = 0;
    assign fifo_intf_81.finish = finish;
    csv_file_dump fifo_csv_dumper_81;
    csv_file_dump cstatus_csv_dumper_81;
    df_fifo_monitor fifo_monitor_81;
    df_fifo_intf fifo_intf_82(clock,reset);
    assign fifo_intf_82.rd_en = AESL_inst_myproject.layer2_out_81_U.if_read & AESL_inst_myproject.layer2_out_81_U.if_empty_n;
    assign fifo_intf_82.wr_en = AESL_inst_myproject.layer2_out_81_U.if_write & AESL_inst_myproject.layer2_out_81_U.if_full_n;
    assign fifo_intf_82.fifo_rd_block = 0;
    assign fifo_intf_82.fifo_wr_block = 0;
    assign fifo_intf_82.finish = finish;
    csv_file_dump fifo_csv_dumper_82;
    csv_file_dump cstatus_csv_dumper_82;
    df_fifo_monitor fifo_monitor_82;
    df_fifo_intf fifo_intf_83(clock,reset);
    assign fifo_intf_83.rd_en = AESL_inst_myproject.layer2_out_82_U.if_read & AESL_inst_myproject.layer2_out_82_U.if_empty_n;
    assign fifo_intf_83.wr_en = AESL_inst_myproject.layer2_out_82_U.if_write & AESL_inst_myproject.layer2_out_82_U.if_full_n;
    assign fifo_intf_83.fifo_rd_block = 0;
    assign fifo_intf_83.fifo_wr_block = 0;
    assign fifo_intf_83.finish = finish;
    csv_file_dump fifo_csv_dumper_83;
    csv_file_dump cstatus_csv_dumper_83;
    df_fifo_monitor fifo_monitor_83;
    df_fifo_intf fifo_intf_84(clock,reset);
    assign fifo_intf_84.rd_en = AESL_inst_myproject.layer2_out_83_U.if_read & AESL_inst_myproject.layer2_out_83_U.if_empty_n;
    assign fifo_intf_84.wr_en = AESL_inst_myproject.layer2_out_83_U.if_write & AESL_inst_myproject.layer2_out_83_U.if_full_n;
    assign fifo_intf_84.fifo_rd_block = 0;
    assign fifo_intf_84.fifo_wr_block = 0;
    assign fifo_intf_84.finish = finish;
    csv_file_dump fifo_csv_dumper_84;
    csv_file_dump cstatus_csv_dumper_84;
    df_fifo_monitor fifo_monitor_84;
    df_fifo_intf fifo_intf_85(clock,reset);
    assign fifo_intf_85.rd_en = AESL_inst_myproject.layer2_out_84_U.if_read & AESL_inst_myproject.layer2_out_84_U.if_empty_n;
    assign fifo_intf_85.wr_en = AESL_inst_myproject.layer2_out_84_U.if_write & AESL_inst_myproject.layer2_out_84_U.if_full_n;
    assign fifo_intf_85.fifo_rd_block = 0;
    assign fifo_intf_85.fifo_wr_block = 0;
    assign fifo_intf_85.finish = finish;
    csv_file_dump fifo_csv_dumper_85;
    csv_file_dump cstatus_csv_dumper_85;
    df_fifo_monitor fifo_monitor_85;
    df_fifo_intf fifo_intf_86(clock,reset);
    assign fifo_intf_86.rd_en = AESL_inst_myproject.layer2_out_85_U.if_read & AESL_inst_myproject.layer2_out_85_U.if_empty_n;
    assign fifo_intf_86.wr_en = AESL_inst_myproject.layer2_out_85_U.if_write & AESL_inst_myproject.layer2_out_85_U.if_full_n;
    assign fifo_intf_86.fifo_rd_block = 0;
    assign fifo_intf_86.fifo_wr_block = 0;
    assign fifo_intf_86.finish = finish;
    csv_file_dump fifo_csv_dumper_86;
    csv_file_dump cstatus_csv_dumper_86;
    df_fifo_monitor fifo_monitor_86;
    df_fifo_intf fifo_intf_87(clock,reset);
    assign fifo_intf_87.rd_en = AESL_inst_myproject.layer2_out_86_U.if_read & AESL_inst_myproject.layer2_out_86_U.if_empty_n;
    assign fifo_intf_87.wr_en = AESL_inst_myproject.layer2_out_86_U.if_write & AESL_inst_myproject.layer2_out_86_U.if_full_n;
    assign fifo_intf_87.fifo_rd_block = 0;
    assign fifo_intf_87.fifo_wr_block = 0;
    assign fifo_intf_87.finish = finish;
    csv_file_dump fifo_csv_dumper_87;
    csv_file_dump cstatus_csv_dumper_87;
    df_fifo_monitor fifo_monitor_87;
    df_fifo_intf fifo_intf_88(clock,reset);
    assign fifo_intf_88.rd_en = AESL_inst_myproject.layer2_out_87_U.if_read & AESL_inst_myproject.layer2_out_87_U.if_empty_n;
    assign fifo_intf_88.wr_en = AESL_inst_myproject.layer2_out_87_U.if_write & AESL_inst_myproject.layer2_out_87_U.if_full_n;
    assign fifo_intf_88.fifo_rd_block = 0;
    assign fifo_intf_88.fifo_wr_block = 0;
    assign fifo_intf_88.finish = finish;
    csv_file_dump fifo_csv_dumper_88;
    csv_file_dump cstatus_csv_dumper_88;
    df_fifo_monitor fifo_monitor_88;
    df_fifo_intf fifo_intf_89(clock,reset);
    assign fifo_intf_89.rd_en = AESL_inst_myproject.layer2_out_88_U.if_read & AESL_inst_myproject.layer2_out_88_U.if_empty_n;
    assign fifo_intf_89.wr_en = AESL_inst_myproject.layer2_out_88_U.if_write & AESL_inst_myproject.layer2_out_88_U.if_full_n;
    assign fifo_intf_89.fifo_rd_block = 0;
    assign fifo_intf_89.fifo_wr_block = 0;
    assign fifo_intf_89.finish = finish;
    csv_file_dump fifo_csv_dumper_89;
    csv_file_dump cstatus_csv_dumper_89;
    df_fifo_monitor fifo_monitor_89;
    df_fifo_intf fifo_intf_90(clock,reset);
    assign fifo_intf_90.rd_en = AESL_inst_myproject.layer2_out_89_U.if_read & AESL_inst_myproject.layer2_out_89_U.if_empty_n;
    assign fifo_intf_90.wr_en = AESL_inst_myproject.layer2_out_89_U.if_write & AESL_inst_myproject.layer2_out_89_U.if_full_n;
    assign fifo_intf_90.fifo_rd_block = 0;
    assign fifo_intf_90.fifo_wr_block = 0;
    assign fifo_intf_90.finish = finish;
    csv_file_dump fifo_csv_dumper_90;
    csv_file_dump cstatus_csv_dumper_90;
    df_fifo_monitor fifo_monitor_90;
    df_fifo_intf fifo_intf_91(clock,reset);
    assign fifo_intf_91.rd_en = AESL_inst_myproject.layer2_out_90_U.if_read & AESL_inst_myproject.layer2_out_90_U.if_empty_n;
    assign fifo_intf_91.wr_en = AESL_inst_myproject.layer2_out_90_U.if_write & AESL_inst_myproject.layer2_out_90_U.if_full_n;
    assign fifo_intf_91.fifo_rd_block = 0;
    assign fifo_intf_91.fifo_wr_block = 0;
    assign fifo_intf_91.finish = finish;
    csv_file_dump fifo_csv_dumper_91;
    csv_file_dump cstatus_csv_dumper_91;
    df_fifo_monitor fifo_monitor_91;
    df_fifo_intf fifo_intf_92(clock,reset);
    assign fifo_intf_92.rd_en = AESL_inst_myproject.layer2_out_91_U.if_read & AESL_inst_myproject.layer2_out_91_U.if_empty_n;
    assign fifo_intf_92.wr_en = AESL_inst_myproject.layer2_out_91_U.if_write & AESL_inst_myproject.layer2_out_91_U.if_full_n;
    assign fifo_intf_92.fifo_rd_block = 0;
    assign fifo_intf_92.fifo_wr_block = 0;
    assign fifo_intf_92.finish = finish;
    csv_file_dump fifo_csv_dumper_92;
    csv_file_dump cstatus_csv_dumper_92;
    df_fifo_monitor fifo_monitor_92;
    df_fifo_intf fifo_intf_93(clock,reset);
    assign fifo_intf_93.rd_en = AESL_inst_myproject.layer2_out_92_U.if_read & AESL_inst_myproject.layer2_out_92_U.if_empty_n;
    assign fifo_intf_93.wr_en = AESL_inst_myproject.layer2_out_92_U.if_write & AESL_inst_myproject.layer2_out_92_U.if_full_n;
    assign fifo_intf_93.fifo_rd_block = 0;
    assign fifo_intf_93.fifo_wr_block = 0;
    assign fifo_intf_93.finish = finish;
    csv_file_dump fifo_csv_dumper_93;
    csv_file_dump cstatus_csv_dumper_93;
    df_fifo_monitor fifo_monitor_93;
    df_fifo_intf fifo_intf_94(clock,reset);
    assign fifo_intf_94.rd_en = AESL_inst_myproject.layer2_out_93_U.if_read & AESL_inst_myproject.layer2_out_93_U.if_empty_n;
    assign fifo_intf_94.wr_en = AESL_inst_myproject.layer2_out_93_U.if_write & AESL_inst_myproject.layer2_out_93_U.if_full_n;
    assign fifo_intf_94.fifo_rd_block = 0;
    assign fifo_intf_94.fifo_wr_block = 0;
    assign fifo_intf_94.finish = finish;
    csv_file_dump fifo_csv_dumper_94;
    csv_file_dump cstatus_csv_dumper_94;
    df_fifo_monitor fifo_monitor_94;
    df_fifo_intf fifo_intf_95(clock,reset);
    assign fifo_intf_95.rd_en = AESL_inst_myproject.layer2_out_94_U.if_read & AESL_inst_myproject.layer2_out_94_U.if_empty_n;
    assign fifo_intf_95.wr_en = AESL_inst_myproject.layer2_out_94_U.if_write & AESL_inst_myproject.layer2_out_94_U.if_full_n;
    assign fifo_intf_95.fifo_rd_block = 0;
    assign fifo_intf_95.fifo_wr_block = 0;
    assign fifo_intf_95.finish = finish;
    csv_file_dump fifo_csv_dumper_95;
    csv_file_dump cstatus_csv_dumper_95;
    df_fifo_monitor fifo_monitor_95;
    df_fifo_intf fifo_intf_96(clock,reset);
    assign fifo_intf_96.rd_en = AESL_inst_myproject.layer2_out_95_U.if_read & AESL_inst_myproject.layer2_out_95_U.if_empty_n;
    assign fifo_intf_96.wr_en = AESL_inst_myproject.layer2_out_95_U.if_write & AESL_inst_myproject.layer2_out_95_U.if_full_n;
    assign fifo_intf_96.fifo_rd_block = 0;
    assign fifo_intf_96.fifo_wr_block = 0;
    assign fifo_intf_96.finish = finish;
    csv_file_dump fifo_csv_dumper_96;
    csv_file_dump cstatus_csv_dumper_96;
    df_fifo_monitor fifo_monitor_96;
    df_fifo_intf fifo_intf_97(clock,reset);
    assign fifo_intf_97.rd_en = AESL_inst_myproject.layer2_out_96_U.if_read & AESL_inst_myproject.layer2_out_96_U.if_empty_n;
    assign fifo_intf_97.wr_en = AESL_inst_myproject.layer2_out_96_U.if_write & AESL_inst_myproject.layer2_out_96_U.if_full_n;
    assign fifo_intf_97.fifo_rd_block = 0;
    assign fifo_intf_97.fifo_wr_block = 0;
    assign fifo_intf_97.finish = finish;
    csv_file_dump fifo_csv_dumper_97;
    csv_file_dump cstatus_csv_dumper_97;
    df_fifo_monitor fifo_monitor_97;
    df_fifo_intf fifo_intf_98(clock,reset);
    assign fifo_intf_98.rd_en = AESL_inst_myproject.layer2_out_97_U.if_read & AESL_inst_myproject.layer2_out_97_U.if_empty_n;
    assign fifo_intf_98.wr_en = AESL_inst_myproject.layer2_out_97_U.if_write & AESL_inst_myproject.layer2_out_97_U.if_full_n;
    assign fifo_intf_98.fifo_rd_block = 0;
    assign fifo_intf_98.fifo_wr_block = 0;
    assign fifo_intf_98.finish = finish;
    csv_file_dump fifo_csv_dumper_98;
    csv_file_dump cstatus_csv_dumper_98;
    df_fifo_monitor fifo_monitor_98;
    df_fifo_intf fifo_intf_99(clock,reset);
    assign fifo_intf_99.rd_en = AESL_inst_myproject.layer2_out_98_U.if_read & AESL_inst_myproject.layer2_out_98_U.if_empty_n;
    assign fifo_intf_99.wr_en = AESL_inst_myproject.layer2_out_98_U.if_write & AESL_inst_myproject.layer2_out_98_U.if_full_n;
    assign fifo_intf_99.fifo_rd_block = 0;
    assign fifo_intf_99.fifo_wr_block = 0;
    assign fifo_intf_99.finish = finish;
    csv_file_dump fifo_csv_dumper_99;
    csv_file_dump cstatus_csv_dumper_99;
    df_fifo_monitor fifo_monitor_99;
    df_fifo_intf fifo_intf_100(clock,reset);
    assign fifo_intf_100.rd_en = AESL_inst_myproject.layer2_out_99_U.if_read & AESL_inst_myproject.layer2_out_99_U.if_empty_n;
    assign fifo_intf_100.wr_en = AESL_inst_myproject.layer2_out_99_U.if_write & AESL_inst_myproject.layer2_out_99_U.if_full_n;
    assign fifo_intf_100.fifo_rd_block = 0;
    assign fifo_intf_100.fifo_wr_block = 0;
    assign fifo_intf_100.finish = finish;
    csv_file_dump fifo_csv_dumper_100;
    csv_file_dump cstatus_csv_dumper_100;
    df_fifo_monitor fifo_monitor_100;
    df_fifo_intf fifo_intf_101(clock,reset);
    assign fifo_intf_101.rd_en = AESL_inst_myproject.layer2_out_100_U.if_read & AESL_inst_myproject.layer2_out_100_U.if_empty_n;
    assign fifo_intf_101.wr_en = AESL_inst_myproject.layer2_out_100_U.if_write & AESL_inst_myproject.layer2_out_100_U.if_full_n;
    assign fifo_intf_101.fifo_rd_block = 0;
    assign fifo_intf_101.fifo_wr_block = 0;
    assign fifo_intf_101.finish = finish;
    csv_file_dump fifo_csv_dumper_101;
    csv_file_dump cstatus_csv_dumper_101;
    df_fifo_monitor fifo_monitor_101;
    df_fifo_intf fifo_intf_102(clock,reset);
    assign fifo_intf_102.rd_en = AESL_inst_myproject.layer2_out_101_U.if_read & AESL_inst_myproject.layer2_out_101_U.if_empty_n;
    assign fifo_intf_102.wr_en = AESL_inst_myproject.layer2_out_101_U.if_write & AESL_inst_myproject.layer2_out_101_U.if_full_n;
    assign fifo_intf_102.fifo_rd_block = 0;
    assign fifo_intf_102.fifo_wr_block = 0;
    assign fifo_intf_102.finish = finish;
    csv_file_dump fifo_csv_dumper_102;
    csv_file_dump cstatus_csv_dumper_102;
    df_fifo_monitor fifo_monitor_102;
    df_fifo_intf fifo_intf_103(clock,reset);
    assign fifo_intf_103.rd_en = AESL_inst_myproject.layer2_out_102_U.if_read & AESL_inst_myproject.layer2_out_102_U.if_empty_n;
    assign fifo_intf_103.wr_en = AESL_inst_myproject.layer2_out_102_U.if_write & AESL_inst_myproject.layer2_out_102_U.if_full_n;
    assign fifo_intf_103.fifo_rd_block = 0;
    assign fifo_intf_103.fifo_wr_block = 0;
    assign fifo_intf_103.finish = finish;
    csv_file_dump fifo_csv_dumper_103;
    csv_file_dump cstatus_csv_dumper_103;
    df_fifo_monitor fifo_monitor_103;
    df_fifo_intf fifo_intf_104(clock,reset);
    assign fifo_intf_104.rd_en = AESL_inst_myproject.layer2_out_103_U.if_read & AESL_inst_myproject.layer2_out_103_U.if_empty_n;
    assign fifo_intf_104.wr_en = AESL_inst_myproject.layer2_out_103_U.if_write & AESL_inst_myproject.layer2_out_103_U.if_full_n;
    assign fifo_intf_104.fifo_rd_block = 0;
    assign fifo_intf_104.fifo_wr_block = 0;
    assign fifo_intf_104.finish = finish;
    csv_file_dump fifo_csv_dumper_104;
    csv_file_dump cstatus_csv_dumper_104;
    df_fifo_monitor fifo_monitor_104;
    df_fifo_intf fifo_intf_105(clock,reset);
    assign fifo_intf_105.rd_en = AESL_inst_myproject.layer2_out_104_U.if_read & AESL_inst_myproject.layer2_out_104_U.if_empty_n;
    assign fifo_intf_105.wr_en = AESL_inst_myproject.layer2_out_104_U.if_write & AESL_inst_myproject.layer2_out_104_U.if_full_n;
    assign fifo_intf_105.fifo_rd_block = 0;
    assign fifo_intf_105.fifo_wr_block = 0;
    assign fifo_intf_105.finish = finish;
    csv_file_dump fifo_csv_dumper_105;
    csv_file_dump cstatus_csv_dumper_105;
    df_fifo_monitor fifo_monitor_105;
    df_fifo_intf fifo_intf_106(clock,reset);
    assign fifo_intf_106.rd_en = AESL_inst_myproject.layer2_out_105_U.if_read & AESL_inst_myproject.layer2_out_105_U.if_empty_n;
    assign fifo_intf_106.wr_en = AESL_inst_myproject.layer2_out_105_U.if_write & AESL_inst_myproject.layer2_out_105_U.if_full_n;
    assign fifo_intf_106.fifo_rd_block = 0;
    assign fifo_intf_106.fifo_wr_block = 0;
    assign fifo_intf_106.finish = finish;
    csv_file_dump fifo_csv_dumper_106;
    csv_file_dump cstatus_csv_dumper_106;
    df_fifo_monitor fifo_monitor_106;
    df_fifo_intf fifo_intf_107(clock,reset);
    assign fifo_intf_107.rd_en = AESL_inst_myproject.layer2_out_106_U.if_read & AESL_inst_myproject.layer2_out_106_U.if_empty_n;
    assign fifo_intf_107.wr_en = AESL_inst_myproject.layer2_out_106_U.if_write & AESL_inst_myproject.layer2_out_106_U.if_full_n;
    assign fifo_intf_107.fifo_rd_block = 0;
    assign fifo_intf_107.fifo_wr_block = 0;
    assign fifo_intf_107.finish = finish;
    csv_file_dump fifo_csv_dumper_107;
    csv_file_dump cstatus_csv_dumper_107;
    df_fifo_monitor fifo_monitor_107;
    df_fifo_intf fifo_intf_108(clock,reset);
    assign fifo_intf_108.rd_en = AESL_inst_myproject.layer2_out_107_U.if_read & AESL_inst_myproject.layer2_out_107_U.if_empty_n;
    assign fifo_intf_108.wr_en = AESL_inst_myproject.layer2_out_107_U.if_write & AESL_inst_myproject.layer2_out_107_U.if_full_n;
    assign fifo_intf_108.fifo_rd_block = 0;
    assign fifo_intf_108.fifo_wr_block = 0;
    assign fifo_intf_108.finish = finish;
    csv_file_dump fifo_csv_dumper_108;
    csv_file_dump cstatus_csv_dumper_108;
    df_fifo_monitor fifo_monitor_108;
    df_fifo_intf fifo_intf_109(clock,reset);
    assign fifo_intf_109.rd_en = AESL_inst_myproject.layer2_out_108_U.if_read & AESL_inst_myproject.layer2_out_108_U.if_empty_n;
    assign fifo_intf_109.wr_en = AESL_inst_myproject.layer2_out_108_U.if_write & AESL_inst_myproject.layer2_out_108_U.if_full_n;
    assign fifo_intf_109.fifo_rd_block = 0;
    assign fifo_intf_109.fifo_wr_block = 0;
    assign fifo_intf_109.finish = finish;
    csv_file_dump fifo_csv_dumper_109;
    csv_file_dump cstatus_csv_dumper_109;
    df_fifo_monitor fifo_monitor_109;
    df_fifo_intf fifo_intf_110(clock,reset);
    assign fifo_intf_110.rd_en = AESL_inst_myproject.layer2_out_109_U.if_read & AESL_inst_myproject.layer2_out_109_U.if_empty_n;
    assign fifo_intf_110.wr_en = AESL_inst_myproject.layer2_out_109_U.if_write & AESL_inst_myproject.layer2_out_109_U.if_full_n;
    assign fifo_intf_110.fifo_rd_block = 0;
    assign fifo_intf_110.fifo_wr_block = 0;
    assign fifo_intf_110.finish = finish;
    csv_file_dump fifo_csv_dumper_110;
    csv_file_dump cstatus_csv_dumper_110;
    df_fifo_monitor fifo_monitor_110;
    df_fifo_intf fifo_intf_111(clock,reset);
    assign fifo_intf_111.rd_en = AESL_inst_myproject.layer2_out_110_U.if_read & AESL_inst_myproject.layer2_out_110_U.if_empty_n;
    assign fifo_intf_111.wr_en = AESL_inst_myproject.layer2_out_110_U.if_write & AESL_inst_myproject.layer2_out_110_U.if_full_n;
    assign fifo_intf_111.fifo_rd_block = 0;
    assign fifo_intf_111.fifo_wr_block = 0;
    assign fifo_intf_111.finish = finish;
    csv_file_dump fifo_csv_dumper_111;
    csv_file_dump cstatus_csv_dumper_111;
    df_fifo_monitor fifo_monitor_111;
    df_fifo_intf fifo_intf_112(clock,reset);
    assign fifo_intf_112.rd_en = AESL_inst_myproject.layer2_out_111_U.if_read & AESL_inst_myproject.layer2_out_111_U.if_empty_n;
    assign fifo_intf_112.wr_en = AESL_inst_myproject.layer2_out_111_U.if_write & AESL_inst_myproject.layer2_out_111_U.if_full_n;
    assign fifo_intf_112.fifo_rd_block = 0;
    assign fifo_intf_112.fifo_wr_block = 0;
    assign fifo_intf_112.finish = finish;
    csv_file_dump fifo_csv_dumper_112;
    csv_file_dump cstatus_csv_dumper_112;
    df_fifo_monitor fifo_monitor_112;
    df_fifo_intf fifo_intf_113(clock,reset);
    assign fifo_intf_113.rd_en = AESL_inst_myproject.layer2_out_112_U.if_read & AESL_inst_myproject.layer2_out_112_U.if_empty_n;
    assign fifo_intf_113.wr_en = AESL_inst_myproject.layer2_out_112_U.if_write & AESL_inst_myproject.layer2_out_112_U.if_full_n;
    assign fifo_intf_113.fifo_rd_block = 0;
    assign fifo_intf_113.fifo_wr_block = 0;
    assign fifo_intf_113.finish = finish;
    csv_file_dump fifo_csv_dumper_113;
    csv_file_dump cstatus_csv_dumper_113;
    df_fifo_monitor fifo_monitor_113;
    df_fifo_intf fifo_intf_114(clock,reset);
    assign fifo_intf_114.rd_en = AESL_inst_myproject.layer2_out_113_U.if_read & AESL_inst_myproject.layer2_out_113_U.if_empty_n;
    assign fifo_intf_114.wr_en = AESL_inst_myproject.layer2_out_113_U.if_write & AESL_inst_myproject.layer2_out_113_U.if_full_n;
    assign fifo_intf_114.fifo_rd_block = 0;
    assign fifo_intf_114.fifo_wr_block = 0;
    assign fifo_intf_114.finish = finish;
    csv_file_dump fifo_csv_dumper_114;
    csv_file_dump cstatus_csv_dumper_114;
    df_fifo_monitor fifo_monitor_114;
    df_fifo_intf fifo_intf_115(clock,reset);
    assign fifo_intf_115.rd_en = AESL_inst_myproject.layer2_out_114_U.if_read & AESL_inst_myproject.layer2_out_114_U.if_empty_n;
    assign fifo_intf_115.wr_en = AESL_inst_myproject.layer2_out_114_U.if_write & AESL_inst_myproject.layer2_out_114_U.if_full_n;
    assign fifo_intf_115.fifo_rd_block = 0;
    assign fifo_intf_115.fifo_wr_block = 0;
    assign fifo_intf_115.finish = finish;
    csv_file_dump fifo_csv_dumper_115;
    csv_file_dump cstatus_csv_dumper_115;
    df_fifo_monitor fifo_monitor_115;
    df_fifo_intf fifo_intf_116(clock,reset);
    assign fifo_intf_116.rd_en = AESL_inst_myproject.layer2_out_115_U.if_read & AESL_inst_myproject.layer2_out_115_U.if_empty_n;
    assign fifo_intf_116.wr_en = AESL_inst_myproject.layer2_out_115_U.if_write & AESL_inst_myproject.layer2_out_115_U.if_full_n;
    assign fifo_intf_116.fifo_rd_block = 0;
    assign fifo_intf_116.fifo_wr_block = 0;
    assign fifo_intf_116.finish = finish;
    csv_file_dump fifo_csv_dumper_116;
    csv_file_dump cstatus_csv_dumper_116;
    df_fifo_monitor fifo_monitor_116;
    df_fifo_intf fifo_intf_117(clock,reset);
    assign fifo_intf_117.rd_en = AESL_inst_myproject.layer2_out_116_U.if_read & AESL_inst_myproject.layer2_out_116_U.if_empty_n;
    assign fifo_intf_117.wr_en = AESL_inst_myproject.layer2_out_116_U.if_write & AESL_inst_myproject.layer2_out_116_U.if_full_n;
    assign fifo_intf_117.fifo_rd_block = 0;
    assign fifo_intf_117.fifo_wr_block = 0;
    assign fifo_intf_117.finish = finish;
    csv_file_dump fifo_csv_dumper_117;
    csv_file_dump cstatus_csv_dumper_117;
    df_fifo_monitor fifo_monitor_117;
    df_fifo_intf fifo_intf_118(clock,reset);
    assign fifo_intf_118.rd_en = AESL_inst_myproject.layer2_out_117_U.if_read & AESL_inst_myproject.layer2_out_117_U.if_empty_n;
    assign fifo_intf_118.wr_en = AESL_inst_myproject.layer2_out_117_U.if_write & AESL_inst_myproject.layer2_out_117_U.if_full_n;
    assign fifo_intf_118.fifo_rd_block = 0;
    assign fifo_intf_118.fifo_wr_block = 0;
    assign fifo_intf_118.finish = finish;
    csv_file_dump fifo_csv_dumper_118;
    csv_file_dump cstatus_csv_dumper_118;
    df_fifo_monitor fifo_monitor_118;
    df_fifo_intf fifo_intf_119(clock,reset);
    assign fifo_intf_119.rd_en = AESL_inst_myproject.layer2_out_118_U.if_read & AESL_inst_myproject.layer2_out_118_U.if_empty_n;
    assign fifo_intf_119.wr_en = AESL_inst_myproject.layer2_out_118_U.if_write & AESL_inst_myproject.layer2_out_118_U.if_full_n;
    assign fifo_intf_119.fifo_rd_block = 0;
    assign fifo_intf_119.fifo_wr_block = 0;
    assign fifo_intf_119.finish = finish;
    csv_file_dump fifo_csv_dumper_119;
    csv_file_dump cstatus_csv_dumper_119;
    df_fifo_monitor fifo_monitor_119;
    df_fifo_intf fifo_intf_120(clock,reset);
    assign fifo_intf_120.rd_en = AESL_inst_myproject.layer2_out_119_U.if_read & AESL_inst_myproject.layer2_out_119_U.if_empty_n;
    assign fifo_intf_120.wr_en = AESL_inst_myproject.layer2_out_119_U.if_write & AESL_inst_myproject.layer2_out_119_U.if_full_n;
    assign fifo_intf_120.fifo_rd_block = 0;
    assign fifo_intf_120.fifo_wr_block = 0;
    assign fifo_intf_120.finish = finish;
    csv_file_dump fifo_csv_dumper_120;
    csv_file_dump cstatus_csv_dumper_120;
    df_fifo_monitor fifo_monitor_120;
    df_fifo_intf fifo_intf_121(clock,reset);
    assign fifo_intf_121.rd_en = AESL_inst_myproject.layer2_out_120_U.if_read & AESL_inst_myproject.layer2_out_120_U.if_empty_n;
    assign fifo_intf_121.wr_en = AESL_inst_myproject.layer2_out_120_U.if_write & AESL_inst_myproject.layer2_out_120_U.if_full_n;
    assign fifo_intf_121.fifo_rd_block = 0;
    assign fifo_intf_121.fifo_wr_block = 0;
    assign fifo_intf_121.finish = finish;
    csv_file_dump fifo_csv_dumper_121;
    csv_file_dump cstatus_csv_dumper_121;
    df_fifo_monitor fifo_monitor_121;
    df_fifo_intf fifo_intf_122(clock,reset);
    assign fifo_intf_122.rd_en = AESL_inst_myproject.layer2_out_121_U.if_read & AESL_inst_myproject.layer2_out_121_U.if_empty_n;
    assign fifo_intf_122.wr_en = AESL_inst_myproject.layer2_out_121_U.if_write & AESL_inst_myproject.layer2_out_121_U.if_full_n;
    assign fifo_intf_122.fifo_rd_block = 0;
    assign fifo_intf_122.fifo_wr_block = 0;
    assign fifo_intf_122.finish = finish;
    csv_file_dump fifo_csv_dumper_122;
    csv_file_dump cstatus_csv_dumper_122;
    df_fifo_monitor fifo_monitor_122;
    df_fifo_intf fifo_intf_123(clock,reset);
    assign fifo_intf_123.rd_en = AESL_inst_myproject.layer2_out_122_U.if_read & AESL_inst_myproject.layer2_out_122_U.if_empty_n;
    assign fifo_intf_123.wr_en = AESL_inst_myproject.layer2_out_122_U.if_write & AESL_inst_myproject.layer2_out_122_U.if_full_n;
    assign fifo_intf_123.fifo_rd_block = 0;
    assign fifo_intf_123.fifo_wr_block = 0;
    assign fifo_intf_123.finish = finish;
    csv_file_dump fifo_csv_dumper_123;
    csv_file_dump cstatus_csv_dumper_123;
    df_fifo_monitor fifo_monitor_123;
    df_fifo_intf fifo_intf_124(clock,reset);
    assign fifo_intf_124.rd_en = AESL_inst_myproject.layer2_out_123_U.if_read & AESL_inst_myproject.layer2_out_123_U.if_empty_n;
    assign fifo_intf_124.wr_en = AESL_inst_myproject.layer2_out_123_U.if_write & AESL_inst_myproject.layer2_out_123_U.if_full_n;
    assign fifo_intf_124.fifo_rd_block = 0;
    assign fifo_intf_124.fifo_wr_block = 0;
    assign fifo_intf_124.finish = finish;
    csv_file_dump fifo_csv_dumper_124;
    csv_file_dump cstatus_csv_dumper_124;
    df_fifo_monitor fifo_monitor_124;
    df_fifo_intf fifo_intf_125(clock,reset);
    assign fifo_intf_125.rd_en = AESL_inst_myproject.layer2_out_124_U.if_read & AESL_inst_myproject.layer2_out_124_U.if_empty_n;
    assign fifo_intf_125.wr_en = AESL_inst_myproject.layer2_out_124_U.if_write & AESL_inst_myproject.layer2_out_124_U.if_full_n;
    assign fifo_intf_125.fifo_rd_block = 0;
    assign fifo_intf_125.fifo_wr_block = 0;
    assign fifo_intf_125.finish = finish;
    csv_file_dump fifo_csv_dumper_125;
    csv_file_dump cstatus_csv_dumper_125;
    df_fifo_monitor fifo_monitor_125;
    df_fifo_intf fifo_intf_126(clock,reset);
    assign fifo_intf_126.rd_en = AESL_inst_myproject.layer2_out_125_U.if_read & AESL_inst_myproject.layer2_out_125_U.if_empty_n;
    assign fifo_intf_126.wr_en = AESL_inst_myproject.layer2_out_125_U.if_write & AESL_inst_myproject.layer2_out_125_U.if_full_n;
    assign fifo_intf_126.fifo_rd_block = 0;
    assign fifo_intf_126.fifo_wr_block = 0;
    assign fifo_intf_126.finish = finish;
    csv_file_dump fifo_csv_dumper_126;
    csv_file_dump cstatus_csv_dumper_126;
    df_fifo_monitor fifo_monitor_126;
    df_fifo_intf fifo_intf_127(clock,reset);
    assign fifo_intf_127.rd_en = AESL_inst_myproject.layer2_out_126_U.if_read & AESL_inst_myproject.layer2_out_126_U.if_empty_n;
    assign fifo_intf_127.wr_en = AESL_inst_myproject.layer2_out_126_U.if_write & AESL_inst_myproject.layer2_out_126_U.if_full_n;
    assign fifo_intf_127.fifo_rd_block = 0;
    assign fifo_intf_127.fifo_wr_block = 0;
    assign fifo_intf_127.finish = finish;
    csv_file_dump fifo_csv_dumper_127;
    csv_file_dump cstatus_csv_dumper_127;
    df_fifo_monitor fifo_monitor_127;
    df_fifo_intf fifo_intf_128(clock,reset);
    assign fifo_intf_128.rd_en = AESL_inst_myproject.layer2_out_127_U.if_read & AESL_inst_myproject.layer2_out_127_U.if_empty_n;
    assign fifo_intf_128.wr_en = AESL_inst_myproject.layer2_out_127_U.if_write & AESL_inst_myproject.layer2_out_127_U.if_full_n;
    assign fifo_intf_128.fifo_rd_block = 0;
    assign fifo_intf_128.fifo_wr_block = 0;
    assign fifo_intf_128.finish = finish;
    csv_file_dump fifo_csv_dumper_128;
    csv_file_dump cstatus_csv_dumper_128;
    df_fifo_monitor fifo_monitor_128;
    df_fifo_intf fifo_intf_129(clock,reset);
    assign fifo_intf_129.rd_en = AESL_inst_myproject.layer2_out_128_U.if_read & AESL_inst_myproject.layer2_out_128_U.if_empty_n;
    assign fifo_intf_129.wr_en = AESL_inst_myproject.layer2_out_128_U.if_write & AESL_inst_myproject.layer2_out_128_U.if_full_n;
    assign fifo_intf_129.fifo_rd_block = 0;
    assign fifo_intf_129.fifo_wr_block = 0;
    assign fifo_intf_129.finish = finish;
    csv_file_dump fifo_csv_dumper_129;
    csv_file_dump cstatus_csv_dumper_129;
    df_fifo_monitor fifo_monitor_129;
    df_fifo_intf fifo_intf_130(clock,reset);
    assign fifo_intf_130.rd_en = AESL_inst_myproject.layer2_out_129_U.if_read & AESL_inst_myproject.layer2_out_129_U.if_empty_n;
    assign fifo_intf_130.wr_en = AESL_inst_myproject.layer2_out_129_U.if_write & AESL_inst_myproject.layer2_out_129_U.if_full_n;
    assign fifo_intf_130.fifo_rd_block = 0;
    assign fifo_intf_130.fifo_wr_block = 0;
    assign fifo_intf_130.finish = finish;
    csv_file_dump fifo_csv_dumper_130;
    csv_file_dump cstatus_csv_dumper_130;
    df_fifo_monitor fifo_monitor_130;
    df_fifo_intf fifo_intf_131(clock,reset);
    assign fifo_intf_131.rd_en = AESL_inst_myproject.layer2_out_130_U.if_read & AESL_inst_myproject.layer2_out_130_U.if_empty_n;
    assign fifo_intf_131.wr_en = AESL_inst_myproject.layer2_out_130_U.if_write & AESL_inst_myproject.layer2_out_130_U.if_full_n;
    assign fifo_intf_131.fifo_rd_block = 0;
    assign fifo_intf_131.fifo_wr_block = 0;
    assign fifo_intf_131.finish = finish;
    csv_file_dump fifo_csv_dumper_131;
    csv_file_dump cstatus_csv_dumper_131;
    df_fifo_monitor fifo_monitor_131;
    df_fifo_intf fifo_intf_132(clock,reset);
    assign fifo_intf_132.rd_en = AESL_inst_myproject.layer2_out_131_U.if_read & AESL_inst_myproject.layer2_out_131_U.if_empty_n;
    assign fifo_intf_132.wr_en = AESL_inst_myproject.layer2_out_131_U.if_write & AESL_inst_myproject.layer2_out_131_U.if_full_n;
    assign fifo_intf_132.fifo_rd_block = 0;
    assign fifo_intf_132.fifo_wr_block = 0;
    assign fifo_intf_132.finish = finish;
    csv_file_dump fifo_csv_dumper_132;
    csv_file_dump cstatus_csv_dumper_132;
    df_fifo_monitor fifo_monitor_132;
    df_fifo_intf fifo_intf_133(clock,reset);
    assign fifo_intf_133.rd_en = AESL_inst_myproject.layer2_out_132_U.if_read & AESL_inst_myproject.layer2_out_132_U.if_empty_n;
    assign fifo_intf_133.wr_en = AESL_inst_myproject.layer2_out_132_U.if_write & AESL_inst_myproject.layer2_out_132_U.if_full_n;
    assign fifo_intf_133.fifo_rd_block = 0;
    assign fifo_intf_133.fifo_wr_block = 0;
    assign fifo_intf_133.finish = finish;
    csv_file_dump fifo_csv_dumper_133;
    csv_file_dump cstatus_csv_dumper_133;
    df_fifo_monitor fifo_monitor_133;
    df_fifo_intf fifo_intf_134(clock,reset);
    assign fifo_intf_134.rd_en = AESL_inst_myproject.layer2_out_133_U.if_read & AESL_inst_myproject.layer2_out_133_U.if_empty_n;
    assign fifo_intf_134.wr_en = AESL_inst_myproject.layer2_out_133_U.if_write & AESL_inst_myproject.layer2_out_133_U.if_full_n;
    assign fifo_intf_134.fifo_rd_block = 0;
    assign fifo_intf_134.fifo_wr_block = 0;
    assign fifo_intf_134.finish = finish;
    csv_file_dump fifo_csv_dumper_134;
    csv_file_dump cstatus_csv_dumper_134;
    df_fifo_monitor fifo_monitor_134;
    df_fifo_intf fifo_intf_135(clock,reset);
    assign fifo_intf_135.rd_en = AESL_inst_myproject.layer2_out_134_U.if_read & AESL_inst_myproject.layer2_out_134_U.if_empty_n;
    assign fifo_intf_135.wr_en = AESL_inst_myproject.layer2_out_134_U.if_write & AESL_inst_myproject.layer2_out_134_U.if_full_n;
    assign fifo_intf_135.fifo_rd_block = 0;
    assign fifo_intf_135.fifo_wr_block = 0;
    assign fifo_intf_135.finish = finish;
    csv_file_dump fifo_csv_dumper_135;
    csv_file_dump cstatus_csv_dumper_135;
    df_fifo_monitor fifo_monitor_135;
    df_fifo_intf fifo_intf_136(clock,reset);
    assign fifo_intf_136.rd_en = AESL_inst_myproject.layer2_out_135_U.if_read & AESL_inst_myproject.layer2_out_135_U.if_empty_n;
    assign fifo_intf_136.wr_en = AESL_inst_myproject.layer2_out_135_U.if_write & AESL_inst_myproject.layer2_out_135_U.if_full_n;
    assign fifo_intf_136.fifo_rd_block = 0;
    assign fifo_intf_136.fifo_wr_block = 0;
    assign fifo_intf_136.finish = finish;
    csv_file_dump fifo_csv_dumper_136;
    csv_file_dump cstatus_csv_dumper_136;
    df_fifo_monitor fifo_monitor_136;
    df_fifo_intf fifo_intf_137(clock,reset);
    assign fifo_intf_137.rd_en = AESL_inst_myproject.layer2_out_136_U.if_read & AESL_inst_myproject.layer2_out_136_U.if_empty_n;
    assign fifo_intf_137.wr_en = AESL_inst_myproject.layer2_out_136_U.if_write & AESL_inst_myproject.layer2_out_136_U.if_full_n;
    assign fifo_intf_137.fifo_rd_block = 0;
    assign fifo_intf_137.fifo_wr_block = 0;
    assign fifo_intf_137.finish = finish;
    csv_file_dump fifo_csv_dumper_137;
    csv_file_dump cstatus_csv_dumper_137;
    df_fifo_monitor fifo_monitor_137;
    df_fifo_intf fifo_intf_138(clock,reset);
    assign fifo_intf_138.rd_en = AESL_inst_myproject.layer2_out_137_U.if_read & AESL_inst_myproject.layer2_out_137_U.if_empty_n;
    assign fifo_intf_138.wr_en = AESL_inst_myproject.layer2_out_137_U.if_write & AESL_inst_myproject.layer2_out_137_U.if_full_n;
    assign fifo_intf_138.fifo_rd_block = 0;
    assign fifo_intf_138.fifo_wr_block = 0;
    assign fifo_intf_138.finish = finish;
    csv_file_dump fifo_csv_dumper_138;
    csv_file_dump cstatus_csv_dumper_138;
    df_fifo_monitor fifo_monitor_138;
    df_fifo_intf fifo_intf_139(clock,reset);
    assign fifo_intf_139.rd_en = AESL_inst_myproject.layer2_out_138_U.if_read & AESL_inst_myproject.layer2_out_138_U.if_empty_n;
    assign fifo_intf_139.wr_en = AESL_inst_myproject.layer2_out_138_U.if_write & AESL_inst_myproject.layer2_out_138_U.if_full_n;
    assign fifo_intf_139.fifo_rd_block = 0;
    assign fifo_intf_139.fifo_wr_block = 0;
    assign fifo_intf_139.finish = finish;
    csv_file_dump fifo_csv_dumper_139;
    csv_file_dump cstatus_csv_dumper_139;
    df_fifo_monitor fifo_monitor_139;
    df_fifo_intf fifo_intf_140(clock,reset);
    assign fifo_intf_140.rd_en = AESL_inst_myproject.layer2_out_139_U.if_read & AESL_inst_myproject.layer2_out_139_U.if_empty_n;
    assign fifo_intf_140.wr_en = AESL_inst_myproject.layer2_out_139_U.if_write & AESL_inst_myproject.layer2_out_139_U.if_full_n;
    assign fifo_intf_140.fifo_rd_block = 0;
    assign fifo_intf_140.fifo_wr_block = 0;
    assign fifo_intf_140.finish = finish;
    csv_file_dump fifo_csv_dumper_140;
    csv_file_dump cstatus_csv_dumper_140;
    df_fifo_monitor fifo_monitor_140;
    df_fifo_intf fifo_intf_141(clock,reset);
    assign fifo_intf_141.rd_en = AESL_inst_myproject.layer2_out_140_U.if_read & AESL_inst_myproject.layer2_out_140_U.if_empty_n;
    assign fifo_intf_141.wr_en = AESL_inst_myproject.layer2_out_140_U.if_write & AESL_inst_myproject.layer2_out_140_U.if_full_n;
    assign fifo_intf_141.fifo_rd_block = 0;
    assign fifo_intf_141.fifo_wr_block = 0;
    assign fifo_intf_141.finish = finish;
    csv_file_dump fifo_csv_dumper_141;
    csv_file_dump cstatus_csv_dumper_141;
    df_fifo_monitor fifo_monitor_141;
    df_fifo_intf fifo_intf_142(clock,reset);
    assign fifo_intf_142.rd_en = AESL_inst_myproject.layer2_out_141_U.if_read & AESL_inst_myproject.layer2_out_141_U.if_empty_n;
    assign fifo_intf_142.wr_en = AESL_inst_myproject.layer2_out_141_U.if_write & AESL_inst_myproject.layer2_out_141_U.if_full_n;
    assign fifo_intf_142.fifo_rd_block = 0;
    assign fifo_intf_142.fifo_wr_block = 0;
    assign fifo_intf_142.finish = finish;
    csv_file_dump fifo_csv_dumper_142;
    csv_file_dump cstatus_csv_dumper_142;
    df_fifo_monitor fifo_monitor_142;
    df_fifo_intf fifo_intf_143(clock,reset);
    assign fifo_intf_143.rd_en = AESL_inst_myproject.layer2_out_142_U.if_read & AESL_inst_myproject.layer2_out_142_U.if_empty_n;
    assign fifo_intf_143.wr_en = AESL_inst_myproject.layer2_out_142_U.if_write & AESL_inst_myproject.layer2_out_142_U.if_full_n;
    assign fifo_intf_143.fifo_rd_block = 0;
    assign fifo_intf_143.fifo_wr_block = 0;
    assign fifo_intf_143.finish = finish;
    csv_file_dump fifo_csv_dumper_143;
    csv_file_dump cstatus_csv_dumper_143;
    df_fifo_monitor fifo_monitor_143;
    df_fifo_intf fifo_intf_144(clock,reset);
    assign fifo_intf_144.rd_en = AESL_inst_myproject.layer2_out_143_U.if_read & AESL_inst_myproject.layer2_out_143_U.if_empty_n;
    assign fifo_intf_144.wr_en = AESL_inst_myproject.layer2_out_143_U.if_write & AESL_inst_myproject.layer2_out_143_U.if_full_n;
    assign fifo_intf_144.fifo_rd_block = 0;
    assign fifo_intf_144.fifo_wr_block = 0;
    assign fifo_intf_144.finish = finish;
    csv_file_dump fifo_csv_dumper_144;
    csv_file_dump cstatus_csv_dumper_144;
    df_fifo_monitor fifo_monitor_144;
    df_fifo_intf fifo_intf_145(clock,reset);
    assign fifo_intf_145.rd_en = AESL_inst_myproject.layer2_out_144_U.if_read & AESL_inst_myproject.layer2_out_144_U.if_empty_n;
    assign fifo_intf_145.wr_en = AESL_inst_myproject.layer2_out_144_U.if_write & AESL_inst_myproject.layer2_out_144_U.if_full_n;
    assign fifo_intf_145.fifo_rd_block = 0;
    assign fifo_intf_145.fifo_wr_block = 0;
    assign fifo_intf_145.finish = finish;
    csv_file_dump fifo_csv_dumper_145;
    csv_file_dump cstatus_csv_dumper_145;
    df_fifo_monitor fifo_monitor_145;
    df_fifo_intf fifo_intf_146(clock,reset);
    assign fifo_intf_146.rd_en = AESL_inst_myproject.layer2_out_145_U.if_read & AESL_inst_myproject.layer2_out_145_U.if_empty_n;
    assign fifo_intf_146.wr_en = AESL_inst_myproject.layer2_out_145_U.if_write & AESL_inst_myproject.layer2_out_145_U.if_full_n;
    assign fifo_intf_146.fifo_rd_block = 0;
    assign fifo_intf_146.fifo_wr_block = 0;
    assign fifo_intf_146.finish = finish;
    csv_file_dump fifo_csv_dumper_146;
    csv_file_dump cstatus_csv_dumper_146;
    df_fifo_monitor fifo_monitor_146;
    df_fifo_intf fifo_intf_147(clock,reset);
    assign fifo_intf_147.rd_en = AESL_inst_myproject.layer2_out_146_U.if_read & AESL_inst_myproject.layer2_out_146_U.if_empty_n;
    assign fifo_intf_147.wr_en = AESL_inst_myproject.layer2_out_146_U.if_write & AESL_inst_myproject.layer2_out_146_U.if_full_n;
    assign fifo_intf_147.fifo_rd_block = 0;
    assign fifo_intf_147.fifo_wr_block = 0;
    assign fifo_intf_147.finish = finish;
    csv_file_dump fifo_csv_dumper_147;
    csv_file_dump cstatus_csv_dumper_147;
    df_fifo_monitor fifo_monitor_147;
    df_fifo_intf fifo_intf_148(clock,reset);
    assign fifo_intf_148.rd_en = AESL_inst_myproject.layer2_out_147_U.if_read & AESL_inst_myproject.layer2_out_147_U.if_empty_n;
    assign fifo_intf_148.wr_en = AESL_inst_myproject.layer2_out_147_U.if_write & AESL_inst_myproject.layer2_out_147_U.if_full_n;
    assign fifo_intf_148.fifo_rd_block = 0;
    assign fifo_intf_148.fifo_wr_block = 0;
    assign fifo_intf_148.finish = finish;
    csv_file_dump fifo_csv_dumper_148;
    csv_file_dump cstatus_csv_dumper_148;
    df_fifo_monitor fifo_monitor_148;
    df_fifo_intf fifo_intf_149(clock,reset);
    assign fifo_intf_149.rd_en = AESL_inst_myproject.layer2_out_148_U.if_read & AESL_inst_myproject.layer2_out_148_U.if_empty_n;
    assign fifo_intf_149.wr_en = AESL_inst_myproject.layer2_out_148_U.if_write & AESL_inst_myproject.layer2_out_148_U.if_full_n;
    assign fifo_intf_149.fifo_rd_block = 0;
    assign fifo_intf_149.fifo_wr_block = 0;
    assign fifo_intf_149.finish = finish;
    csv_file_dump fifo_csv_dumper_149;
    csv_file_dump cstatus_csv_dumper_149;
    df_fifo_monitor fifo_monitor_149;
    df_fifo_intf fifo_intf_150(clock,reset);
    assign fifo_intf_150.rd_en = AESL_inst_myproject.layer2_out_149_U.if_read & AESL_inst_myproject.layer2_out_149_U.if_empty_n;
    assign fifo_intf_150.wr_en = AESL_inst_myproject.layer2_out_149_U.if_write & AESL_inst_myproject.layer2_out_149_U.if_full_n;
    assign fifo_intf_150.fifo_rd_block = 0;
    assign fifo_intf_150.fifo_wr_block = 0;
    assign fifo_intf_150.finish = finish;
    csv_file_dump fifo_csv_dumper_150;
    csv_file_dump cstatus_csv_dumper_150;
    df_fifo_monitor fifo_monitor_150;
    df_fifo_intf fifo_intf_151(clock,reset);
    assign fifo_intf_151.rd_en = AESL_inst_myproject.layer2_out_150_U.if_read & AESL_inst_myproject.layer2_out_150_U.if_empty_n;
    assign fifo_intf_151.wr_en = AESL_inst_myproject.layer2_out_150_U.if_write & AESL_inst_myproject.layer2_out_150_U.if_full_n;
    assign fifo_intf_151.fifo_rd_block = 0;
    assign fifo_intf_151.fifo_wr_block = 0;
    assign fifo_intf_151.finish = finish;
    csv_file_dump fifo_csv_dumper_151;
    csv_file_dump cstatus_csv_dumper_151;
    df_fifo_monitor fifo_monitor_151;
    df_fifo_intf fifo_intf_152(clock,reset);
    assign fifo_intf_152.rd_en = AESL_inst_myproject.layer2_out_151_U.if_read & AESL_inst_myproject.layer2_out_151_U.if_empty_n;
    assign fifo_intf_152.wr_en = AESL_inst_myproject.layer2_out_151_U.if_write & AESL_inst_myproject.layer2_out_151_U.if_full_n;
    assign fifo_intf_152.fifo_rd_block = 0;
    assign fifo_intf_152.fifo_wr_block = 0;
    assign fifo_intf_152.finish = finish;
    csv_file_dump fifo_csv_dumper_152;
    csv_file_dump cstatus_csv_dumper_152;
    df_fifo_monitor fifo_monitor_152;
    df_fifo_intf fifo_intf_153(clock,reset);
    assign fifo_intf_153.rd_en = AESL_inst_myproject.layer2_out_152_U.if_read & AESL_inst_myproject.layer2_out_152_U.if_empty_n;
    assign fifo_intf_153.wr_en = AESL_inst_myproject.layer2_out_152_U.if_write & AESL_inst_myproject.layer2_out_152_U.if_full_n;
    assign fifo_intf_153.fifo_rd_block = 0;
    assign fifo_intf_153.fifo_wr_block = 0;
    assign fifo_intf_153.finish = finish;
    csv_file_dump fifo_csv_dumper_153;
    csv_file_dump cstatus_csv_dumper_153;
    df_fifo_monitor fifo_monitor_153;
    df_fifo_intf fifo_intf_154(clock,reset);
    assign fifo_intf_154.rd_en = AESL_inst_myproject.layer2_out_153_U.if_read & AESL_inst_myproject.layer2_out_153_U.if_empty_n;
    assign fifo_intf_154.wr_en = AESL_inst_myproject.layer2_out_153_U.if_write & AESL_inst_myproject.layer2_out_153_U.if_full_n;
    assign fifo_intf_154.fifo_rd_block = 0;
    assign fifo_intf_154.fifo_wr_block = 0;
    assign fifo_intf_154.finish = finish;
    csv_file_dump fifo_csv_dumper_154;
    csv_file_dump cstatus_csv_dumper_154;
    df_fifo_monitor fifo_monitor_154;
    df_fifo_intf fifo_intf_155(clock,reset);
    assign fifo_intf_155.rd_en = AESL_inst_myproject.layer2_out_154_U.if_read & AESL_inst_myproject.layer2_out_154_U.if_empty_n;
    assign fifo_intf_155.wr_en = AESL_inst_myproject.layer2_out_154_U.if_write & AESL_inst_myproject.layer2_out_154_U.if_full_n;
    assign fifo_intf_155.fifo_rd_block = 0;
    assign fifo_intf_155.fifo_wr_block = 0;
    assign fifo_intf_155.finish = finish;
    csv_file_dump fifo_csv_dumper_155;
    csv_file_dump cstatus_csv_dumper_155;
    df_fifo_monitor fifo_monitor_155;
    df_fifo_intf fifo_intf_156(clock,reset);
    assign fifo_intf_156.rd_en = AESL_inst_myproject.layer2_out_155_U.if_read & AESL_inst_myproject.layer2_out_155_U.if_empty_n;
    assign fifo_intf_156.wr_en = AESL_inst_myproject.layer2_out_155_U.if_write & AESL_inst_myproject.layer2_out_155_U.if_full_n;
    assign fifo_intf_156.fifo_rd_block = 0;
    assign fifo_intf_156.fifo_wr_block = 0;
    assign fifo_intf_156.finish = finish;
    csv_file_dump fifo_csv_dumper_156;
    csv_file_dump cstatus_csv_dumper_156;
    df_fifo_monitor fifo_monitor_156;
    df_fifo_intf fifo_intf_157(clock,reset);
    assign fifo_intf_157.rd_en = AESL_inst_myproject.layer2_out_156_U.if_read & AESL_inst_myproject.layer2_out_156_U.if_empty_n;
    assign fifo_intf_157.wr_en = AESL_inst_myproject.layer2_out_156_U.if_write & AESL_inst_myproject.layer2_out_156_U.if_full_n;
    assign fifo_intf_157.fifo_rd_block = 0;
    assign fifo_intf_157.fifo_wr_block = 0;
    assign fifo_intf_157.finish = finish;
    csv_file_dump fifo_csv_dumper_157;
    csv_file_dump cstatus_csv_dumper_157;
    df_fifo_monitor fifo_monitor_157;
    df_fifo_intf fifo_intf_158(clock,reset);
    assign fifo_intf_158.rd_en = AESL_inst_myproject.layer2_out_157_U.if_read & AESL_inst_myproject.layer2_out_157_U.if_empty_n;
    assign fifo_intf_158.wr_en = AESL_inst_myproject.layer2_out_157_U.if_write & AESL_inst_myproject.layer2_out_157_U.if_full_n;
    assign fifo_intf_158.fifo_rd_block = 0;
    assign fifo_intf_158.fifo_wr_block = 0;
    assign fifo_intf_158.finish = finish;
    csv_file_dump fifo_csv_dumper_158;
    csv_file_dump cstatus_csv_dumper_158;
    df_fifo_monitor fifo_monitor_158;
    df_fifo_intf fifo_intf_159(clock,reset);
    assign fifo_intf_159.rd_en = AESL_inst_myproject.layer2_out_158_U.if_read & AESL_inst_myproject.layer2_out_158_U.if_empty_n;
    assign fifo_intf_159.wr_en = AESL_inst_myproject.layer2_out_158_U.if_write & AESL_inst_myproject.layer2_out_158_U.if_full_n;
    assign fifo_intf_159.fifo_rd_block = 0;
    assign fifo_intf_159.fifo_wr_block = 0;
    assign fifo_intf_159.finish = finish;
    csv_file_dump fifo_csv_dumper_159;
    csv_file_dump cstatus_csv_dumper_159;
    df_fifo_monitor fifo_monitor_159;
    df_fifo_intf fifo_intf_160(clock,reset);
    assign fifo_intf_160.rd_en = AESL_inst_myproject.layer2_out_159_U.if_read & AESL_inst_myproject.layer2_out_159_U.if_empty_n;
    assign fifo_intf_160.wr_en = AESL_inst_myproject.layer2_out_159_U.if_write & AESL_inst_myproject.layer2_out_159_U.if_full_n;
    assign fifo_intf_160.fifo_rd_block = 0;
    assign fifo_intf_160.fifo_wr_block = 0;
    assign fifo_intf_160.finish = finish;
    csv_file_dump fifo_csv_dumper_160;
    csv_file_dump cstatus_csv_dumper_160;
    df_fifo_monitor fifo_monitor_160;
    df_fifo_intf fifo_intf_161(clock,reset);
    assign fifo_intf_161.rd_en = AESL_inst_myproject.layer2_out_160_U.if_read & AESL_inst_myproject.layer2_out_160_U.if_empty_n;
    assign fifo_intf_161.wr_en = AESL_inst_myproject.layer2_out_160_U.if_write & AESL_inst_myproject.layer2_out_160_U.if_full_n;
    assign fifo_intf_161.fifo_rd_block = 0;
    assign fifo_intf_161.fifo_wr_block = 0;
    assign fifo_intf_161.finish = finish;
    csv_file_dump fifo_csv_dumper_161;
    csv_file_dump cstatus_csv_dumper_161;
    df_fifo_monitor fifo_monitor_161;
    df_fifo_intf fifo_intf_162(clock,reset);
    assign fifo_intf_162.rd_en = AESL_inst_myproject.layer2_out_161_U.if_read & AESL_inst_myproject.layer2_out_161_U.if_empty_n;
    assign fifo_intf_162.wr_en = AESL_inst_myproject.layer2_out_161_U.if_write & AESL_inst_myproject.layer2_out_161_U.if_full_n;
    assign fifo_intf_162.fifo_rd_block = 0;
    assign fifo_intf_162.fifo_wr_block = 0;
    assign fifo_intf_162.finish = finish;
    csv_file_dump fifo_csv_dumper_162;
    csv_file_dump cstatus_csv_dumper_162;
    df_fifo_monitor fifo_monitor_162;
    df_fifo_intf fifo_intf_163(clock,reset);
    assign fifo_intf_163.rd_en = AESL_inst_myproject.layer2_out_162_U.if_read & AESL_inst_myproject.layer2_out_162_U.if_empty_n;
    assign fifo_intf_163.wr_en = AESL_inst_myproject.layer2_out_162_U.if_write & AESL_inst_myproject.layer2_out_162_U.if_full_n;
    assign fifo_intf_163.fifo_rd_block = 0;
    assign fifo_intf_163.fifo_wr_block = 0;
    assign fifo_intf_163.finish = finish;
    csv_file_dump fifo_csv_dumper_163;
    csv_file_dump cstatus_csv_dumper_163;
    df_fifo_monitor fifo_monitor_163;
    df_fifo_intf fifo_intf_164(clock,reset);
    assign fifo_intf_164.rd_en = AESL_inst_myproject.layer2_out_163_U.if_read & AESL_inst_myproject.layer2_out_163_U.if_empty_n;
    assign fifo_intf_164.wr_en = AESL_inst_myproject.layer2_out_163_U.if_write & AESL_inst_myproject.layer2_out_163_U.if_full_n;
    assign fifo_intf_164.fifo_rd_block = 0;
    assign fifo_intf_164.fifo_wr_block = 0;
    assign fifo_intf_164.finish = finish;
    csv_file_dump fifo_csv_dumper_164;
    csv_file_dump cstatus_csv_dumper_164;
    df_fifo_monitor fifo_monitor_164;
    df_fifo_intf fifo_intf_165(clock,reset);
    assign fifo_intf_165.rd_en = AESL_inst_myproject.layer2_out_164_U.if_read & AESL_inst_myproject.layer2_out_164_U.if_empty_n;
    assign fifo_intf_165.wr_en = AESL_inst_myproject.layer2_out_164_U.if_write & AESL_inst_myproject.layer2_out_164_U.if_full_n;
    assign fifo_intf_165.fifo_rd_block = 0;
    assign fifo_intf_165.fifo_wr_block = 0;
    assign fifo_intf_165.finish = finish;
    csv_file_dump fifo_csv_dumper_165;
    csv_file_dump cstatus_csv_dumper_165;
    df_fifo_monitor fifo_monitor_165;
    df_fifo_intf fifo_intf_166(clock,reset);
    assign fifo_intf_166.rd_en = AESL_inst_myproject.layer2_out_165_U.if_read & AESL_inst_myproject.layer2_out_165_U.if_empty_n;
    assign fifo_intf_166.wr_en = AESL_inst_myproject.layer2_out_165_U.if_write & AESL_inst_myproject.layer2_out_165_U.if_full_n;
    assign fifo_intf_166.fifo_rd_block = 0;
    assign fifo_intf_166.fifo_wr_block = 0;
    assign fifo_intf_166.finish = finish;
    csv_file_dump fifo_csv_dumper_166;
    csv_file_dump cstatus_csv_dumper_166;
    df_fifo_monitor fifo_monitor_166;
    df_fifo_intf fifo_intf_167(clock,reset);
    assign fifo_intf_167.rd_en = AESL_inst_myproject.layer2_out_166_U.if_read & AESL_inst_myproject.layer2_out_166_U.if_empty_n;
    assign fifo_intf_167.wr_en = AESL_inst_myproject.layer2_out_166_U.if_write & AESL_inst_myproject.layer2_out_166_U.if_full_n;
    assign fifo_intf_167.fifo_rd_block = 0;
    assign fifo_intf_167.fifo_wr_block = 0;
    assign fifo_intf_167.finish = finish;
    csv_file_dump fifo_csv_dumper_167;
    csv_file_dump cstatus_csv_dumper_167;
    df_fifo_monitor fifo_monitor_167;
    df_fifo_intf fifo_intf_168(clock,reset);
    assign fifo_intf_168.rd_en = AESL_inst_myproject.layer2_out_167_U.if_read & AESL_inst_myproject.layer2_out_167_U.if_empty_n;
    assign fifo_intf_168.wr_en = AESL_inst_myproject.layer2_out_167_U.if_write & AESL_inst_myproject.layer2_out_167_U.if_full_n;
    assign fifo_intf_168.fifo_rd_block = 0;
    assign fifo_intf_168.fifo_wr_block = 0;
    assign fifo_intf_168.finish = finish;
    csv_file_dump fifo_csv_dumper_168;
    csv_file_dump cstatus_csv_dumper_168;
    df_fifo_monitor fifo_monitor_168;
    df_fifo_intf fifo_intf_169(clock,reset);
    assign fifo_intf_169.rd_en = AESL_inst_myproject.layer2_out_168_U.if_read & AESL_inst_myproject.layer2_out_168_U.if_empty_n;
    assign fifo_intf_169.wr_en = AESL_inst_myproject.layer2_out_168_U.if_write & AESL_inst_myproject.layer2_out_168_U.if_full_n;
    assign fifo_intf_169.fifo_rd_block = 0;
    assign fifo_intf_169.fifo_wr_block = 0;
    assign fifo_intf_169.finish = finish;
    csv_file_dump fifo_csv_dumper_169;
    csv_file_dump cstatus_csv_dumper_169;
    df_fifo_monitor fifo_monitor_169;
    df_fifo_intf fifo_intf_170(clock,reset);
    assign fifo_intf_170.rd_en = AESL_inst_myproject.layer2_out_169_U.if_read & AESL_inst_myproject.layer2_out_169_U.if_empty_n;
    assign fifo_intf_170.wr_en = AESL_inst_myproject.layer2_out_169_U.if_write & AESL_inst_myproject.layer2_out_169_U.if_full_n;
    assign fifo_intf_170.fifo_rd_block = 0;
    assign fifo_intf_170.fifo_wr_block = 0;
    assign fifo_intf_170.finish = finish;
    csv_file_dump fifo_csv_dumper_170;
    csv_file_dump cstatus_csv_dumper_170;
    df_fifo_monitor fifo_monitor_170;
    df_fifo_intf fifo_intf_171(clock,reset);
    assign fifo_intf_171.rd_en = AESL_inst_myproject.layer2_out_170_U.if_read & AESL_inst_myproject.layer2_out_170_U.if_empty_n;
    assign fifo_intf_171.wr_en = AESL_inst_myproject.layer2_out_170_U.if_write & AESL_inst_myproject.layer2_out_170_U.if_full_n;
    assign fifo_intf_171.fifo_rd_block = 0;
    assign fifo_intf_171.fifo_wr_block = 0;
    assign fifo_intf_171.finish = finish;
    csv_file_dump fifo_csv_dumper_171;
    csv_file_dump cstatus_csv_dumper_171;
    df_fifo_monitor fifo_monitor_171;
    df_fifo_intf fifo_intf_172(clock,reset);
    assign fifo_intf_172.rd_en = AESL_inst_myproject.layer2_out_171_U.if_read & AESL_inst_myproject.layer2_out_171_U.if_empty_n;
    assign fifo_intf_172.wr_en = AESL_inst_myproject.layer2_out_171_U.if_write & AESL_inst_myproject.layer2_out_171_U.if_full_n;
    assign fifo_intf_172.fifo_rd_block = 0;
    assign fifo_intf_172.fifo_wr_block = 0;
    assign fifo_intf_172.finish = finish;
    csv_file_dump fifo_csv_dumper_172;
    csv_file_dump cstatus_csv_dumper_172;
    df_fifo_monitor fifo_monitor_172;
    df_fifo_intf fifo_intf_173(clock,reset);
    assign fifo_intf_173.rd_en = AESL_inst_myproject.layer2_out_172_U.if_read & AESL_inst_myproject.layer2_out_172_U.if_empty_n;
    assign fifo_intf_173.wr_en = AESL_inst_myproject.layer2_out_172_U.if_write & AESL_inst_myproject.layer2_out_172_U.if_full_n;
    assign fifo_intf_173.fifo_rd_block = 0;
    assign fifo_intf_173.fifo_wr_block = 0;
    assign fifo_intf_173.finish = finish;
    csv_file_dump fifo_csv_dumper_173;
    csv_file_dump cstatus_csv_dumper_173;
    df_fifo_monitor fifo_monitor_173;
    df_fifo_intf fifo_intf_174(clock,reset);
    assign fifo_intf_174.rd_en = AESL_inst_myproject.layer2_out_173_U.if_read & AESL_inst_myproject.layer2_out_173_U.if_empty_n;
    assign fifo_intf_174.wr_en = AESL_inst_myproject.layer2_out_173_U.if_write & AESL_inst_myproject.layer2_out_173_U.if_full_n;
    assign fifo_intf_174.fifo_rd_block = 0;
    assign fifo_intf_174.fifo_wr_block = 0;
    assign fifo_intf_174.finish = finish;
    csv_file_dump fifo_csv_dumper_174;
    csv_file_dump cstatus_csv_dumper_174;
    df_fifo_monitor fifo_monitor_174;
    df_fifo_intf fifo_intf_175(clock,reset);
    assign fifo_intf_175.rd_en = AESL_inst_myproject.layer2_out_174_U.if_read & AESL_inst_myproject.layer2_out_174_U.if_empty_n;
    assign fifo_intf_175.wr_en = AESL_inst_myproject.layer2_out_174_U.if_write & AESL_inst_myproject.layer2_out_174_U.if_full_n;
    assign fifo_intf_175.fifo_rd_block = 0;
    assign fifo_intf_175.fifo_wr_block = 0;
    assign fifo_intf_175.finish = finish;
    csv_file_dump fifo_csv_dumper_175;
    csv_file_dump cstatus_csv_dumper_175;
    df_fifo_monitor fifo_monitor_175;
    df_fifo_intf fifo_intf_176(clock,reset);
    assign fifo_intf_176.rd_en = AESL_inst_myproject.layer2_out_175_U.if_read & AESL_inst_myproject.layer2_out_175_U.if_empty_n;
    assign fifo_intf_176.wr_en = AESL_inst_myproject.layer2_out_175_U.if_write & AESL_inst_myproject.layer2_out_175_U.if_full_n;
    assign fifo_intf_176.fifo_rd_block = 0;
    assign fifo_intf_176.fifo_wr_block = 0;
    assign fifo_intf_176.finish = finish;
    csv_file_dump fifo_csv_dumper_176;
    csv_file_dump cstatus_csv_dumper_176;
    df_fifo_monitor fifo_monitor_176;
    df_fifo_intf fifo_intf_177(clock,reset);
    assign fifo_intf_177.rd_en = AESL_inst_myproject.layer2_out_176_U.if_read & AESL_inst_myproject.layer2_out_176_U.if_empty_n;
    assign fifo_intf_177.wr_en = AESL_inst_myproject.layer2_out_176_U.if_write & AESL_inst_myproject.layer2_out_176_U.if_full_n;
    assign fifo_intf_177.fifo_rd_block = 0;
    assign fifo_intf_177.fifo_wr_block = 0;
    assign fifo_intf_177.finish = finish;
    csv_file_dump fifo_csv_dumper_177;
    csv_file_dump cstatus_csv_dumper_177;
    df_fifo_monitor fifo_monitor_177;
    df_fifo_intf fifo_intf_178(clock,reset);
    assign fifo_intf_178.rd_en = AESL_inst_myproject.layer2_out_177_U.if_read & AESL_inst_myproject.layer2_out_177_U.if_empty_n;
    assign fifo_intf_178.wr_en = AESL_inst_myproject.layer2_out_177_U.if_write & AESL_inst_myproject.layer2_out_177_U.if_full_n;
    assign fifo_intf_178.fifo_rd_block = 0;
    assign fifo_intf_178.fifo_wr_block = 0;
    assign fifo_intf_178.finish = finish;
    csv_file_dump fifo_csv_dumper_178;
    csv_file_dump cstatus_csv_dumper_178;
    df_fifo_monitor fifo_monitor_178;
    df_fifo_intf fifo_intf_179(clock,reset);
    assign fifo_intf_179.rd_en = AESL_inst_myproject.layer2_out_178_U.if_read & AESL_inst_myproject.layer2_out_178_U.if_empty_n;
    assign fifo_intf_179.wr_en = AESL_inst_myproject.layer2_out_178_U.if_write & AESL_inst_myproject.layer2_out_178_U.if_full_n;
    assign fifo_intf_179.fifo_rd_block = 0;
    assign fifo_intf_179.fifo_wr_block = 0;
    assign fifo_intf_179.finish = finish;
    csv_file_dump fifo_csv_dumper_179;
    csv_file_dump cstatus_csv_dumper_179;
    df_fifo_monitor fifo_monitor_179;
    df_fifo_intf fifo_intf_180(clock,reset);
    assign fifo_intf_180.rd_en = AESL_inst_myproject.layer2_out_179_U.if_read & AESL_inst_myproject.layer2_out_179_U.if_empty_n;
    assign fifo_intf_180.wr_en = AESL_inst_myproject.layer2_out_179_U.if_write & AESL_inst_myproject.layer2_out_179_U.if_full_n;
    assign fifo_intf_180.fifo_rd_block = 0;
    assign fifo_intf_180.fifo_wr_block = 0;
    assign fifo_intf_180.finish = finish;
    csv_file_dump fifo_csv_dumper_180;
    csv_file_dump cstatus_csv_dumper_180;
    df_fifo_monitor fifo_monitor_180;
    df_fifo_intf fifo_intf_181(clock,reset);
    assign fifo_intf_181.rd_en = AESL_inst_myproject.layer2_out_180_U.if_read & AESL_inst_myproject.layer2_out_180_U.if_empty_n;
    assign fifo_intf_181.wr_en = AESL_inst_myproject.layer2_out_180_U.if_write & AESL_inst_myproject.layer2_out_180_U.if_full_n;
    assign fifo_intf_181.fifo_rd_block = 0;
    assign fifo_intf_181.fifo_wr_block = 0;
    assign fifo_intf_181.finish = finish;
    csv_file_dump fifo_csv_dumper_181;
    csv_file_dump cstatus_csv_dumper_181;
    df_fifo_monitor fifo_monitor_181;
    df_fifo_intf fifo_intf_182(clock,reset);
    assign fifo_intf_182.rd_en = AESL_inst_myproject.layer2_out_181_U.if_read & AESL_inst_myproject.layer2_out_181_U.if_empty_n;
    assign fifo_intf_182.wr_en = AESL_inst_myproject.layer2_out_181_U.if_write & AESL_inst_myproject.layer2_out_181_U.if_full_n;
    assign fifo_intf_182.fifo_rd_block = 0;
    assign fifo_intf_182.fifo_wr_block = 0;
    assign fifo_intf_182.finish = finish;
    csv_file_dump fifo_csv_dumper_182;
    csv_file_dump cstatus_csv_dumper_182;
    df_fifo_monitor fifo_monitor_182;
    df_fifo_intf fifo_intf_183(clock,reset);
    assign fifo_intf_183.rd_en = AESL_inst_myproject.layer2_out_182_U.if_read & AESL_inst_myproject.layer2_out_182_U.if_empty_n;
    assign fifo_intf_183.wr_en = AESL_inst_myproject.layer2_out_182_U.if_write & AESL_inst_myproject.layer2_out_182_U.if_full_n;
    assign fifo_intf_183.fifo_rd_block = 0;
    assign fifo_intf_183.fifo_wr_block = 0;
    assign fifo_intf_183.finish = finish;
    csv_file_dump fifo_csv_dumper_183;
    csv_file_dump cstatus_csv_dumper_183;
    df_fifo_monitor fifo_monitor_183;
    df_fifo_intf fifo_intf_184(clock,reset);
    assign fifo_intf_184.rd_en = AESL_inst_myproject.layer2_out_183_U.if_read & AESL_inst_myproject.layer2_out_183_U.if_empty_n;
    assign fifo_intf_184.wr_en = AESL_inst_myproject.layer2_out_183_U.if_write & AESL_inst_myproject.layer2_out_183_U.if_full_n;
    assign fifo_intf_184.fifo_rd_block = 0;
    assign fifo_intf_184.fifo_wr_block = 0;
    assign fifo_intf_184.finish = finish;
    csv_file_dump fifo_csv_dumper_184;
    csv_file_dump cstatus_csv_dumper_184;
    df_fifo_monitor fifo_monitor_184;
    df_fifo_intf fifo_intf_185(clock,reset);
    assign fifo_intf_185.rd_en = AESL_inst_myproject.layer2_out_184_U.if_read & AESL_inst_myproject.layer2_out_184_U.if_empty_n;
    assign fifo_intf_185.wr_en = AESL_inst_myproject.layer2_out_184_U.if_write & AESL_inst_myproject.layer2_out_184_U.if_full_n;
    assign fifo_intf_185.fifo_rd_block = 0;
    assign fifo_intf_185.fifo_wr_block = 0;
    assign fifo_intf_185.finish = finish;
    csv_file_dump fifo_csv_dumper_185;
    csv_file_dump cstatus_csv_dumper_185;
    df_fifo_monitor fifo_monitor_185;
    df_fifo_intf fifo_intf_186(clock,reset);
    assign fifo_intf_186.rd_en = AESL_inst_myproject.layer2_out_185_U.if_read & AESL_inst_myproject.layer2_out_185_U.if_empty_n;
    assign fifo_intf_186.wr_en = AESL_inst_myproject.layer2_out_185_U.if_write & AESL_inst_myproject.layer2_out_185_U.if_full_n;
    assign fifo_intf_186.fifo_rd_block = 0;
    assign fifo_intf_186.fifo_wr_block = 0;
    assign fifo_intf_186.finish = finish;
    csv_file_dump fifo_csv_dumper_186;
    csv_file_dump cstatus_csv_dumper_186;
    df_fifo_monitor fifo_monitor_186;
    df_fifo_intf fifo_intf_187(clock,reset);
    assign fifo_intf_187.rd_en = AESL_inst_myproject.layer2_out_186_U.if_read & AESL_inst_myproject.layer2_out_186_U.if_empty_n;
    assign fifo_intf_187.wr_en = AESL_inst_myproject.layer2_out_186_U.if_write & AESL_inst_myproject.layer2_out_186_U.if_full_n;
    assign fifo_intf_187.fifo_rd_block = 0;
    assign fifo_intf_187.fifo_wr_block = 0;
    assign fifo_intf_187.finish = finish;
    csv_file_dump fifo_csv_dumper_187;
    csv_file_dump cstatus_csv_dumper_187;
    df_fifo_monitor fifo_monitor_187;
    df_fifo_intf fifo_intf_188(clock,reset);
    assign fifo_intf_188.rd_en = AESL_inst_myproject.layer2_out_187_U.if_read & AESL_inst_myproject.layer2_out_187_U.if_empty_n;
    assign fifo_intf_188.wr_en = AESL_inst_myproject.layer2_out_187_U.if_write & AESL_inst_myproject.layer2_out_187_U.if_full_n;
    assign fifo_intf_188.fifo_rd_block = 0;
    assign fifo_intf_188.fifo_wr_block = 0;
    assign fifo_intf_188.finish = finish;
    csv_file_dump fifo_csv_dumper_188;
    csv_file_dump cstatus_csv_dumper_188;
    df_fifo_monitor fifo_monitor_188;
    df_fifo_intf fifo_intf_189(clock,reset);
    assign fifo_intf_189.rd_en = AESL_inst_myproject.layer2_out_188_U.if_read & AESL_inst_myproject.layer2_out_188_U.if_empty_n;
    assign fifo_intf_189.wr_en = AESL_inst_myproject.layer2_out_188_U.if_write & AESL_inst_myproject.layer2_out_188_U.if_full_n;
    assign fifo_intf_189.fifo_rd_block = 0;
    assign fifo_intf_189.fifo_wr_block = 0;
    assign fifo_intf_189.finish = finish;
    csv_file_dump fifo_csv_dumper_189;
    csv_file_dump cstatus_csv_dumper_189;
    df_fifo_monitor fifo_monitor_189;
    df_fifo_intf fifo_intf_190(clock,reset);
    assign fifo_intf_190.rd_en = AESL_inst_myproject.layer2_out_189_U.if_read & AESL_inst_myproject.layer2_out_189_U.if_empty_n;
    assign fifo_intf_190.wr_en = AESL_inst_myproject.layer2_out_189_U.if_write & AESL_inst_myproject.layer2_out_189_U.if_full_n;
    assign fifo_intf_190.fifo_rd_block = 0;
    assign fifo_intf_190.fifo_wr_block = 0;
    assign fifo_intf_190.finish = finish;
    csv_file_dump fifo_csv_dumper_190;
    csv_file_dump cstatus_csv_dumper_190;
    df_fifo_monitor fifo_monitor_190;
    df_fifo_intf fifo_intf_191(clock,reset);
    assign fifo_intf_191.rd_en = AESL_inst_myproject.layer2_out_190_U.if_read & AESL_inst_myproject.layer2_out_190_U.if_empty_n;
    assign fifo_intf_191.wr_en = AESL_inst_myproject.layer2_out_190_U.if_write & AESL_inst_myproject.layer2_out_190_U.if_full_n;
    assign fifo_intf_191.fifo_rd_block = 0;
    assign fifo_intf_191.fifo_wr_block = 0;
    assign fifo_intf_191.finish = finish;
    csv_file_dump fifo_csv_dumper_191;
    csv_file_dump cstatus_csv_dumper_191;
    df_fifo_monitor fifo_monitor_191;
    df_fifo_intf fifo_intf_192(clock,reset);
    assign fifo_intf_192.rd_en = AESL_inst_myproject.layer2_out_191_U.if_read & AESL_inst_myproject.layer2_out_191_U.if_empty_n;
    assign fifo_intf_192.wr_en = AESL_inst_myproject.layer2_out_191_U.if_write & AESL_inst_myproject.layer2_out_191_U.if_full_n;
    assign fifo_intf_192.fifo_rd_block = 0;
    assign fifo_intf_192.fifo_wr_block = 0;
    assign fifo_intf_192.finish = finish;
    csv_file_dump fifo_csv_dumper_192;
    csv_file_dump cstatus_csv_dumper_192;
    df_fifo_monitor fifo_monitor_192;
    df_fifo_intf fifo_intf_193(clock,reset);
    assign fifo_intf_193.rd_en = AESL_inst_myproject.layer2_out_192_U.if_read & AESL_inst_myproject.layer2_out_192_U.if_empty_n;
    assign fifo_intf_193.wr_en = AESL_inst_myproject.layer2_out_192_U.if_write & AESL_inst_myproject.layer2_out_192_U.if_full_n;
    assign fifo_intf_193.fifo_rd_block = 0;
    assign fifo_intf_193.fifo_wr_block = 0;
    assign fifo_intf_193.finish = finish;
    csv_file_dump fifo_csv_dumper_193;
    csv_file_dump cstatus_csv_dumper_193;
    df_fifo_monitor fifo_monitor_193;
    df_fifo_intf fifo_intf_194(clock,reset);
    assign fifo_intf_194.rd_en = AESL_inst_myproject.layer2_out_193_U.if_read & AESL_inst_myproject.layer2_out_193_U.if_empty_n;
    assign fifo_intf_194.wr_en = AESL_inst_myproject.layer2_out_193_U.if_write & AESL_inst_myproject.layer2_out_193_U.if_full_n;
    assign fifo_intf_194.fifo_rd_block = 0;
    assign fifo_intf_194.fifo_wr_block = 0;
    assign fifo_intf_194.finish = finish;
    csv_file_dump fifo_csv_dumper_194;
    csv_file_dump cstatus_csv_dumper_194;
    df_fifo_monitor fifo_monitor_194;
    df_fifo_intf fifo_intf_195(clock,reset);
    assign fifo_intf_195.rd_en = AESL_inst_myproject.layer2_out_194_U.if_read & AESL_inst_myproject.layer2_out_194_U.if_empty_n;
    assign fifo_intf_195.wr_en = AESL_inst_myproject.layer2_out_194_U.if_write & AESL_inst_myproject.layer2_out_194_U.if_full_n;
    assign fifo_intf_195.fifo_rd_block = 0;
    assign fifo_intf_195.fifo_wr_block = 0;
    assign fifo_intf_195.finish = finish;
    csv_file_dump fifo_csv_dumper_195;
    csv_file_dump cstatus_csv_dumper_195;
    df_fifo_monitor fifo_monitor_195;
    df_fifo_intf fifo_intf_196(clock,reset);
    assign fifo_intf_196.rd_en = AESL_inst_myproject.layer2_out_195_U.if_read & AESL_inst_myproject.layer2_out_195_U.if_empty_n;
    assign fifo_intf_196.wr_en = AESL_inst_myproject.layer2_out_195_U.if_write & AESL_inst_myproject.layer2_out_195_U.if_full_n;
    assign fifo_intf_196.fifo_rd_block = 0;
    assign fifo_intf_196.fifo_wr_block = 0;
    assign fifo_intf_196.finish = finish;
    csv_file_dump fifo_csv_dumper_196;
    csv_file_dump cstatus_csv_dumper_196;
    df_fifo_monitor fifo_monitor_196;
    df_fifo_intf fifo_intf_197(clock,reset);
    assign fifo_intf_197.rd_en = AESL_inst_myproject.layer2_out_196_U.if_read & AESL_inst_myproject.layer2_out_196_U.if_empty_n;
    assign fifo_intf_197.wr_en = AESL_inst_myproject.layer2_out_196_U.if_write & AESL_inst_myproject.layer2_out_196_U.if_full_n;
    assign fifo_intf_197.fifo_rd_block = 0;
    assign fifo_intf_197.fifo_wr_block = 0;
    assign fifo_intf_197.finish = finish;
    csv_file_dump fifo_csv_dumper_197;
    csv_file_dump cstatus_csv_dumper_197;
    df_fifo_monitor fifo_monitor_197;
    df_fifo_intf fifo_intf_198(clock,reset);
    assign fifo_intf_198.rd_en = AESL_inst_myproject.layer2_out_197_U.if_read & AESL_inst_myproject.layer2_out_197_U.if_empty_n;
    assign fifo_intf_198.wr_en = AESL_inst_myproject.layer2_out_197_U.if_write & AESL_inst_myproject.layer2_out_197_U.if_full_n;
    assign fifo_intf_198.fifo_rd_block = 0;
    assign fifo_intf_198.fifo_wr_block = 0;
    assign fifo_intf_198.finish = finish;
    csv_file_dump fifo_csv_dumper_198;
    csv_file_dump cstatus_csv_dumper_198;
    df_fifo_monitor fifo_monitor_198;
    df_fifo_intf fifo_intf_199(clock,reset);
    assign fifo_intf_199.rd_en = AESL_inst_myproject.layer2_out_198_U.if_read & AESL_inst_myproject.layer2_out_198_U.if_empty_n;
    assign fifo_intf_199.wr_en = AESL_inst_myproject.layer2_out_198_U.if_write & AESL_inst_myproject.layer2_out_198_U.if_full_n;
    assign fifo_intf_199.fifo_rd_block = 0;
    assign fifo_intf_199.fifo_wr_block = 0;
    assign fifo_intf_199.finish = finish;
    csv_file_dump fifo_csv_dumper_199;
    csv_file_dump cstatus_csv_dumper_199;
    df_fifo_monitor fifo_monitor_199;
    df_fifo_intf fifo_intf_200(clock,reset);
    assign fifo_intf_200.rd_en = AESL_inst_myproject.layer2_out_199_U.if_read & AESL_inst_myproject.layer2_out_199_U.if_empty_n;
    assign fifo_intf_200.wr_en = AESL_inst_myproject.layer2_out_199_U.if_write & AESL_inst_myproject.layer2_out_199_U.if_full_n;
    assign fifo_intf_200.fifo_rd_block = 0;
    assign fifo_intf_200.fifo_wr_block = 0;
    assign fifo_intf_200.finish = finish;
    csv_file_dump fifo_csv_dumper_200;
    csv_file_dump cstatus_csv_dumper_200;
    df_fifo_monitor fifo_monitor_200;
    df_fifo_intf fifo_intf_201(clock,reset);
    assign fifo_intf_201.rd_en = AESL_inst_myproject.layer2_out_200_U.if_read & AESL_inst_myproject.layer2_out_200_U.if_empty_n;
    assign fifo_intf_201.wr_en = AESL_inst_myproject.layer2_out_200_U.if_write & AESL_inst_myproject.layer2_out_200_U.if_full_n;
    assign fifo_intf_201.fifo_rd_block = 0;
    assign fifo_intf_201.fifo_wr_block = 0;
    assign fifo_intf_201.finish = finish;
    csv_file_dump fifo_csv_dumper_201;
    csv_file_dump cstatus_csv_dumper_201;
    df_fifo_monitor fifo_monitor_201;
    df_fifo_intf fifo_intf_202(clock,reset);
    assign fifo_intf_202.rd_en = AESL_inst_myproject.layer2_out_201_U.if_read & AESL_inst_myproject.layer2_out_201_U.if_empty_n;
    assign fifo_intf_202.wr_en = AESL_inst_myproject.layer2_out_201_U.if_write & AESL_inst_myproject.layer2_out_201_U.if_full_n;
    assign fifo_intf_202.fifo_rd_block = 0;
    assign fifo_intf_202.fifo_wr_block = 0;
    assign fifo_intf_202.finish = finish;
    csv_file_dump fifo_csv_dumper_202;
    csv_file_dump cstatus_csv_dumper_202;
    df_fifo_monitor fifo_monitor_202;
    df_fifo_intf fifo_intf_203(clock,reset);
    assign fifo_intf_203.rd_en = AESL_inst_myproject.layer2_out_202_U.if_read & AESL_inst_myproject.layer2_out_202_U.if_empty_n;
    assign fifo_intf_203.wr_en = AESL_inst_myproject.layer2_out_202_U.if_write & AESL_inst_myproject.layer2_out_202_U.if_full_n;
    assign fifo_intf_203.fifo_rd_block = 0;
    assign fifo_intf_203.fifo_wr_block = 0;
    assign fifo_intf_203.finish = finish;
    csv_file_dump fifo_csv_dumper_203;
    csv_file_dump cstatus_csv_dumper_203;
    df_fifo_monitor fifo_monitor_203;
    df_fifo_intf fifo_intf_204(clock,reset);
    assign fifo_intf_204.rd_en = AESL_inst_myproject.layer2_out_203_U.if_read & AESL_inst_myproject.layer2_out_203_U.if_empty_n;
    assign fifo_intf_204.wr_en = AESL_inst_myproject.layer2_out_203_U.if_write & AESL_inst_myproject.layer2_out_203_U.if_full_n;
    assign fifo_intf_204.fifo_rd_block = 0;
    assign fifo_intf_204.fifo_wr_block = 0;
    assign fifo_intf_204.finish = finish;
    csv_file_dump fifo_csv_dumper_204;
    csv_file_dump cstatus_csv_dumper_204;
    df_fifo_monitor fifo_monitor_204;
    df_fifo_intf fifo_intf_205(clock,reset);
    assign fifo_intf_205.rd_en = AESL_inst_myproject.layer2_out_204_U.if_read & AESL_inst_myproject.layer2_out_204_U.if_empty_n;
    assign fifo_intf_205.wr_en = AESL_inst_myproject.layer2_out_204_U.if_write & AESL_inst_myproject.layer2_out_204_U.if_full_n;
    assign fifo_intf_205.fifo_rd_block = 0;
    assign fifo_intf_205.fifo_wr_block = 0;
    assign fifo_intf_205.finish = finish;
    csv_file_dump fifo_csv_dumper_205;
    csv_file_dump cstatus_csv_dumper_205;
    df_fifo_monitor fifo_monitor_205;
    df_fifo_intf fifo_intf_206(clock,reset);
    assign fifo_intf_206.rd_en = AESL_inst_myproject.layer2_out_205_U.if_read & AESL_inst_myproject.layer2_out_205_U.if_empty_n;
    assign fifo_intf_206.wr_en = AESL_inst_myproject.layer2_out_205_U.if_write & AESL_inst_myproject.layer2_out_205_U.if_full_n;
    assign fifo_intf_206.fifo_rd_block = 0;
    assign fifo_intf_206.fifo_wr_block = 0;
    assign fifo_intf_206.finish = finish;
    csv_file_dump fifo_csv_dumper_206;
    csv_file_dump cstatus_csv_dumper_206;
    df_fifo_monitor fifo_monitor_206;
    df_fifo_intf fifo_intf_207(clock,reset);
    assign fifo_intf_207.rd_en = AESL_inst_myproject.layer2_out_206_U.if_read & AESL_inst_myproject.layer2_out_206_U.if_empty_n;
    assign fifo_intf_207.wr_en = AESL_inst_myproject.layer2_out_206_U.if_write & AESL_inst_myproject.layer2_out_206_U.if_full_n;
    assign fifo_intf_207.fifo_rd_block = 0;
    assign fifo_intf_207.fifo_wr_block = 0;
    assign fifo_intf_207.finish = finish;
    csv_file_dump fifo_csv_dumper_207;
    csv_file_dump cstatus_csv_dumper_207;
    df_fifo_monitor fifo_monitor_207;
    df_fifo_intf fifo_intf_208(clock,reset);
    assign fifo_intf_208.rd_en = AESL_inst_myproject.layer2_out_207_U.if_read & AESL_inst_myproject.layer2_out_207_U.if_empty_n;
    assign fifo_intf_208.wr_en = AESL_inst_myproject.layer2_out_207_U.if_write & AESL_inst_myproject.layer2_out_207_U.if_full_n;
    assign fifo_intf_208.fifo_rd_block = 0;
    assign fifo_intf_208.fifo_wr_block = 0;
    assign fifo_intf_208.finish = finish;
    csv_file_dump fifo_csv_dumper_208;
    csv_file_dump cstatus_csv_dumper_208;
    df_fifo_monitor fifo_monitor_208;
    df_fifo_intf fifo_intf_209(clock,reset);
    assign fifo_intf_209.rd_en = AESL_inst_myproject.layer2_out_208_U.if_read & AESL_inst_myproject.layer2_out_208_U.if_empty_n;
    assign fifo_intf_209.wr_en = AESL_inst_myproject.layer2_out_208_U.if_write & AESL_inst_myproject.layer2_out_208_U.if_full_n;
    assign fifo_intf_209.fifo_rd_block = 0;
    assign fifo_intf_209.fifo_wr_block = 0;
    assign fifo_intf_209.finish = finish;
    csv_file_dump fifo_csv_dumper_209;
    csv_file_dump cstatus_csv_dumper_209;
    df_fifo_monitor fifo_monitor_209;
    df_fifo_intf fifo_intf_210(clock,reset);
    assign fifo_intf_210.rd_en = AESL_inst_myproject.layer2_out_209_U.if_read & AESL_inst_myproject.layer2_out_209_U.if_empty_n;
    assign fifo_intf_210.wr_en = AESL_inst_myproject.layer2_out_209_U.if_write & AESL_inst_myproject.layer2_out_209_U.if_full_n;
    assign fifo_intf_210.fifo_rd_block = 0;
    assign fifo_intf_210.fifo_wr_block = 0;
    assign fifo_intf_210.finish = finish;
    csv_file_dump fifo_csv_dumper_210;
    csv_file_dump cstatus_csv_dumper_210;
    df_fifo_monitor fifo_monitor_210;
    df_fifo_intf fifo_intf_211(clock,reset);
    assign fifo_intf_211.rd_en = AESL_inst_myproject.layer2_out_210_U.if_read & AESL_inst_myproject.layer2_out_210_U.if_empty_n;
    assign fifo_intf_211.wr_en = AESL_inst_myproject.layer2_out_210_U.if_write & AESL_inst_myproject.layer2_out_210_U.if_full_n;
    assign fifo_intf_211.fifo_rd_block = 0;
    assign fifo_intf_211.fifo_wr_block = 0;
    assign fifo_intf_211.finish = finish;
    csv_file_dump fifo_csv_dumper_211;
    csv_file_dump cstatus_csv_dumper_211;
    df_fifo_monitor fifo_monitor_211;
    df_fifo_intf fifo_intf_212(clock,reset);
    assign fifo_intf_212.rd_en = AESL_inst_myproject.layer2_out_211_U.if_read & AESL_inst_myproject.layer2_out_211_U.if_empty_n;
    assign fifo_intf_212.wr_en = AESL_inst_myproject.layer2_out_211_U.if_write & AESL_inst_myproject.layer2_out_211_U.if_full_n;
    assign fifo_intf_212.fifo_rd_block = 0;
    assign fifo_intf_212.fifo_wr_block = 0;
    assign fifo_intf_212.finish = finish;
    csv_file_dump fifo_csv_dumper_212;
    csv_file_dump cstatus_csv_dumper_212;
    df_fifo_monitor fifo_monitor_212;
    df_fifo_intf fifo_intf_213(clock,reset);
    assign fifo_intf_213.rd_en = AESL_inst_myproject.layer2_out_212_U.if_read & AESL_inst_myproject.layer2_out_212_U.if_empty_n;
    assign fifo_intf_213.wr_en = AESL_inst_myproject.layer2_out_212_U.if_write & AESL_inst_myproject.layer2_out_212_U.if_full_n;
    assign fifo_intf_213.fifo_rd_block = 0;
    assign fifo_intf_213.fifo_wr_block = 0;
    assign fifo_intf_213.finish = finish;
    csv_file_dump fifo_csv_dumper_213;
    csv_file_dump cstatus_csv_dumper_213;
    df_fifo_monitor fifo_monitor_213;
    df_fifo_intf fifo_intf_214(clock,reset);
    assign fifo_intf_214.rd_en = AESL_inst_myproject.layer2_out_213_U.if_read & AESL_inst_myproject.layer2_out_213_U.if_empty_n;
    assign fifo_intf_214.wr_en = AESL_inst_myproject.layer2_out_213_U.if_write & AESL_inst_myproject.layer2_out_213_U.if_full_n;
    assign fifo_intf_214.fifo_rd_block = 0;
    assign fifo_intf_214.fifo_wr_block = 0;
    assign fifo_intf_214.finish = finish;
    csv_file_dump fifo_csv_dumper_214;
    csv_file_dump cstatus_csv_dumper_214;
    df_fifo_monitor fifo_monitor_214;
    df_fifo_intf fifo_intf_215(clock,reset);
    assign fifo_intf_215.rd_en = AESL_inst_myproject.layer2_out_214_U.if_read & AESL_inst_myproject.layer2_out_214_U.if_empty_n;
    assign fifo_intf_215.wr_en = AESL_inst_myproject.layer2_out_214_U.if_write & AESL_inst_myproject.layer2_out_214_U.if_full_n;
    assign fifo_intf_215.fifo_rd_block = 0;
    assign fifo_intf_215.fifo_wr_block = 0;
    assign fifo_intf_215.finish = finish;
    csv_file_dump fifo_csv_dumper_215;
    csv_file_dump cstatus_csv_dumper_215;
    df_fifo_monitor fifo_monitor_215;
    df_fifo_intf fifo_intf_216(clock,reset);
    assign fifo_intf_216.rd_en = AESL_inst_myproject.layer2_out_215_U.if_read & AESL_inst_myproject.layer2_out_215_U.if_empty_n;
    assign fifo_intf_216.wr_en = AESL_inst_myproject.layer2_out_215_U.if_write & AESL_inst_myproject.layer2_out_215_U.if_full_n;
    assign fifo_intf_216.fifo_rd_block = 0;
    assign fifo_intf_216.fifo_wr_block = 0;
    assign fifo_intf_216.finish = finish;
    csv_file_dump fifo_csv_dumper_216;
    csv_file_dump cstatus_csv_dumper_216;
    df_fifo_monitor fifo_monitor_216;
    df_fifo_intf fifo_intf_217(clock,reset);
    assign fifo_intf_217.rd_en = AESL_inst_myproject.layer2_out_216_U.if_read & AESL_inst_myproject.layer2_out_216_U.if_empty_n;
    assign fifo_intf_217.wr_en = AESL_inst_myproject.layer2_out_216_U.if_write & AESL_inst_myproject.layer2_out_216_U.if_full_n;
    assign fifo_intf_217.fifo_rd_block = 0;
    assign fifo_intf_217.fifo_wr_block = 0;
    assign fifo_intf_217.finish = finish;
    csv_file_dump fifo_csv_dumper_217;
    csv_file_dump cstatus_csv_dumper_217;
    df_fifo_monitor fifo_monitor_217;
    df_fifo_intf fifo_intf_218(clock,reset);
    assign fifo_intf_218.rd_en = AESL_inst_myproject.layer2_out_217_U.if_read & AESL_inst_myproject.layer2_out_217_U.if_empty_n;
    assign fifo_intf_218.wr_en = AESL_inst_myproject.layer2_out_217_U.if_write & AESL_inst_myproject.layer2_out_217_U.if_full_n;
    assign fifo_intf_218.fifo_rd_block = 0;
    assign fifo_intf_218.fifo_wr_block = 0;
    assign fifo_intf_218.finish = finish;
    csv_file_dump fifo_csv_dumper_218;
    csv_file_dump cstatus_csv_dumper_218;
    df_fifo_monitor fifo_monitor_218;
    df_fifo_intf fifo_intf_219(clock,reset);
    assign fifo_intf_219.rd_en = AESL_inst_myproject.layer2_out_218_U.if_read & AESL_inst_myproject.layer2_out_218_U.if_empty_n;
    assign fifo_intf_219.wr_en = AESL_inst_myproject.layer2_out_218_U.if_write & AESL_inst_myproject.layer2_out_218_U.if_full_n;
    assign fifo_intf_219.fifo_rd_block = 0;
    assign fifo_intf_219.fifo_wr_block = 0;
    assign fifo_intf_219.finish = finish;
    csv_file_dump fifo_csv_dumper_219;
    csv_file_dump cstatus_csv_dumper_219;
    df_fifo_monitor fifo_monitor_219;
    df_fifo_intf fifo_intf_220(clock,reset);
    assign fifo_intf_220.rd_en = AESL_inst_myproject.layer2_out_219_U.if_read & AESL_inst_myproject.layer2_out_219_U.if_empty_n;
    assign fifo_intf_220.wr_en = AESL_inst_myproject.layer2_out_219_U.if_write & AESL_inst_myproject.layer2_out_219_U.if_full_n;
    assign fifo_intf_220.fifo_rd_block = 0;
    assign fifo_intf_220.fifo_wr_block = 0;
    assign fifo_intf_220.finish = finish;
    csv_file_dump fifo_csv_dumper_220;
    csv_file_dump cstatus_csv_dumper_220;
    df_fifo_monitor fifo_monitor_220;
    df_fifo_intf fifo_intf_221(clock,reset);
    assign fifo_intf_221.rd_en = AESL_inst_myproject.layer2_out_220_U.if_read & AESL_inst_myproject.layer2_out_220_U.if_empty_n;
    assign fifo_intf_221.wr_en = AESL_inst_myproject.layer2_out_220_U.if_write & AESL_inst_myproject.layer2_out_220_U.if_full_n;
    assign fifo_intf_221.fifo_rd_block = 0;
    assign fifo_intf_221.fifo_wr_block = 0;
    assign fifo_intf_221.finish = finish;
    csv_file_dump fifo_csv_dumper_221;
    csv_file_dump cstatus_csv_dumper_221;
    df_fifo_monitor fifo_monitor_221;
    df_fifo_intf fifo_intf_222(clock,reset);
    assign fifo_intf_222.rd_en = AESL_inst_myproject.layer2_out_221_U.if_read & AESL_inst_myproject.layer2_out_221_U.if_empty_n;
    assign fifo_intf_222.wr_en = AESL_inst_myproject.layer2_out_221_U.if_write & AESL_inst_myproject.layer2_out_221_U.if_full_n;
    assign fifo_intf_222.fifo_rd_block = 0;
    assign fifo_intf_222.fifo_wr_block = 0;
    assign fifo_intf_222.finish = finish;
    csv_file_dump fifo_csv_dumper_222;
    csv_file_dump cstatus_csv_dumper_222;
    df_fifo_monitor fifo_monitor_222;
    df_fifo_intf fifo_intf_223(clock,reset);
    assign fifo_intf_223.rd_en = AESL_inst_myproject.layer2_out_222_U.if_read & AESL_inst_myproject.layer2_out_222_U.if_empty_n;
    assign fifo_intf_223.wr_en = AESL_inst_myproject.layer2_out_222_U.if_write & AESL_inst_myproject.layer2_out_222_U.if_full_n;
    assign fifo_intf_223.fifo_rd_block = 0;
    assign fifo_intf_223.fifo_wr_block = 0;
    assign fifo_intf_223.finish = finish;
    csv_file_dump fifo_csv_dumper_223;
    csv_file_dump cstatus_csv_dumper_223;
    df_fifo_monitor fifo_monitor_223;
    df_fifo_intf fifo_intf_224(clock,reset);
    assign fifo_intf_224.rd_en = AESL_inst_myproject.layer2_out_223_U.if_read & AESL_inst_myproject.layer2_out_223_U.if_empty_n;
    assign fifo_intf_224.wr_en = AESL_inst_myproject.layer2_out_223_U.if_write & AESL_inst_myproject.layer2_out_223_U.if_full_n;
    assign fifo_intf_224.fifo_rd_block = 0;
    assign fifo_intf_224.fifo_wr_block = 0;
    assign fifo_intf_224.finish = finish;
    csv_file_dump fifo_csv_dumper_224;
    csv_file_dump cstatus_csv_dumper_224;
    df_fifo_monitor fifo_monitor_224;
    df_fifo_intf fifo_intf_225(clock,reset);
    assign fifo_intf_225.rd_en = AESL_inst_myproject.layer2_out_224_U.if_read & AESL_inst_myproject.layer2_out_224_U.if_empty_n;
    assign fifo_intf_225.wr_en = AESL_inst_myproject.layer2_out_224_U.if_write & AESL_inst_myproject.layer2_out_224_U.if_full_n;
    assign fifo_intf_225.fifo_rd_block = 0;
    assign fifo_intf_225.fifo_wr_block = 0;
    assign fifo_intf_225.finish = finish;
    csv_file_dump fifo_csv_dumper_225;
    csv_file_dump cstatus_csv_dumper_225;
    df_fifo_monitor fifo_monitor_225;
    df_fifo_intf fifo_intf_226(clock,reset);
    assign fifo_intf_226.rd_en = AESL_inst_myproject.layer2_out_225_U.if_read & AESL_inst_myproject.layer2_out_225_U.if_empty_n;
    assign fifo_intf_226.wr_en = AESL_inst_myproject.layer2_out_225_U.if_write & AESL_inst_myproject.layer2_out_225_U.if_full_n;
    assign fifo_intf_226.fifo_rd_block = 0;
    assign fifo_intf_226.fifo_wr_block = 0;
    assign fifo_intf_226.finish = finish;
    csv_file_dump fifo_csv_dumper_226;
    csv_file_dump cstatus_csv_dumper_226;
    df_fifo_monitor fifo_monitor_226;
    df_fifo_intf fifo_intf_227(clock,reset);
    assign fifo_intf_227.rd_en = AESL_inst_myproject.layer2_out_226_U.if_read & AESL_inst_myproject.layer2_out_226_U.if_empty_n;
    assign fifo_intf_227.wr_en = AESL_inst_myproject.layer2_out_226_U.if_write & AESL_inst_myproject.layer2_out_226_U.if_full_n;
    assign fifo_intf_227.fifo_rd_block = 0;
    assign fifo_intf_227.fifo_wr_block = 0;
    assign fifo_intf_227.finish = finish;
    csv_file_dump fifo_csv_dumper_227;
    csv_file_dump cstatus_csv_dumper_227;
    df_fifo_monitor fifo_monitor_227;
    df_fifo_intf fifo_intf_228(clock,reset);
    assign fifo_intf_228.rd_en = AESL_inst_myproject.layer2_out_227_U.if_read & AESL_inst_myproject.layer2_out_227_U.if_empty_n;
    assign fifo_intf_228.wr_en = AESL_inst_myproject.layer2_out_227_U.if_write & AESL_inst_myproject.layer2_out_227_U.if_full_n;
    assign fifo_intf_228.fifo_rd_block = 0;
    assign fifo_intf_228.fifo_wr_block = 0;
    assign fifo_intf_228.finish = finish;
    csv_file_dump fifo_csv_dumper_228;
    csv_file_dump cstatus_csv_dumper_228;
    df_fifo_monitor fifo_monitor_228;
    df_fifo_intf fifo_intf_229(clock,reset);
    assign fifo_intf_229.rd_en = AESL_inst_myproject.layer2_out_228_U.if_read & AESL_inst_myproject.layer2_out_228_U.if_empty_n;
    assign fifo_intf_229.wr_en = AESL_inst_myproject.layer2_out_228_U.if_write & AESL_inst_myproject.layer2_out_228_U.if_full_n;
    assign fifo_intf_229.fifo_rd_block = 0;
    assign fifo_intf_229.fifo_wr_block = 0;
    assign fifo_intf_229.finish = finish;
    csv_file_dump fifo_csv_dumper_229;
    csv_file_dump cstatus_csv_dumper_229;
    df_fifo_monitor fifo_monitor_229;
    df_fifo_intf fifo_intf_230(clock,reset);
    assign fifo_intf_230.rd_en = AESL_inst_myproject.layer2_out_229_U.if_read & AESL_inst_myproject.layer2_out_229_U.if_empty_n;
    assign fifo_intf_230.wr_en = AESL_inst_myproject.layer2_out_229_U.if_write & AESL_inst_myproject.layer2_out_229_U.if_full_n;
    assign fifo_intf_230.fifo_rd_block = 0;
    assign fifo_intf_230.fifo_wr_block = 0;
    assign fifo_intf_230.finish = finish;
    csv_file_dump fifo_csv_dumper_230;
    csv_file_dump cstatus_csv_dumper_230;
    df_fifo_monitor fifo_monitor_230;
    df_fifo_intf fifo_intf_231(clock,reset);
    assign fifo_intf_231.rd_en = AESL_inst_myproject.layer2_out_230_U.if_read & AESL_inst_myproject.layer2_out_230_U.if_empty_n;
    assign fifo_intf_231.wr_en = AESL_inst_myproject.layer2_out_230_U.if_write & AESL_inst_myproject.layer2_out_230_U.if_full_n;
    assign fifo_intf_231.fifo_rd_block = 0;
    assign fifo_intf_231.fifo_wr_block = 0;
    assign fifo_intf_231.finish = finish;
    csv_file_dump fifo_csv_dumper_231;
    csv_file_dump cstatus_csv_dumper_231;
    df_fifo_monitor fifo_monitor_231;
    df_fifo_intf fifo_intf_232(clock,reset);
    assign fifo_intf_232.rd_en = AESL_inst_myproject.layer2_out_231_U.if_read & AESL_inst_myproject.layer2_out_231_U.if_empty_n;
    assign fifo_intf_232.wr_en = AESL_inst_myproject.layer2_out_231_U.if_write & AESL_inst_myproject.layer2_out_231_U.if_full_n;
    assign fifo_intf_232.fifo_rd_block = 0;
    assign fifo_intf_232.fifo_wr_block = 0;
    assign fifo_intf_232.finish = finish;
    csv_file_dump fifo_csv_dumper_232;
    csv_file_dump cstatus_csv_dumper_232;
    df_fifo_monitor fifo_monitor_232;
    df_fifo_intf fifo_intf_233(clock,reset);
    assign fifo_intf_233.rd_en = AESL_inst_myproject.layer2_out_232_U.if_read & AESL_inst_myproject.layer2_out_232_U.if_empty_n;
    assign fifo_intf_233.wr_en = AESL_inst_myproject.layer2_out_232_U.if_write & AESL_inst_myproject.layer2_out_232_U.if_full_n;
    assign fifo_intf_233.fifo_rd_block = 0;
    assign fifo_intf_233.fifo_wr_block = 0;
    assign fifo_intf_233.finish = finish;
    csv_file_dump fifo_csv_dumper_233;
    csv_file_dump cstatus_csv_dumper_233;
    df_fifo_monitor fifo_monitor_233;
    df_fifo_intf fifo_intf_234(clock,reset);
    assign fifo_intf_234.rd_en = AESL_inst_myproject.layer2_out_233_U.if_read & AESL_inst_myproject.layer2_out_233_U.if_empty_n;
    assign fifo_intf_234.wr_en = AESL_inst_myproject.layer2_out_233_U.if_write & AESL_inst_myproject.layer2_out_233_U.if_full_n;
    assign fifo_intf_234.fifo_rd_block = 0;
    assign fifo_intf_234.fifo_wr_block = 0;
    assign fifo_intf_234.finish = finish;
    csv_file_dump fifo_csv_dumper_234;
    csv_file_dump cstatus_csv_dumper_234;
    df_fifo_monitor fifo_monitor_234;
    df_fifo_intf fifo_intf_235(clock,reset);
    assign fifo_intf_235.rd_en = AESL_inst_myproject.layer2_out_234_U.if_read & AESL_inst_myproject.layer2_out_234_U.if_empty_n;
    assign fifo_intf_235.wr_en = AESL_inst_myproject.layer2_out_234_U.if_write & AESL_inst_myproject.layer2_out_234_U.if_full_n;
    assign fifo_intf_235.fifo_rd_block = 0;
    assign fifo_intf_235.fifo_wr_block = 0;
    assign fifo_intf_235.finish = finish;
    csv_file_dump fifo_csv_dumper_235;
    csv_file_dump cstatus_csv_dumper_235;
    df_fifo_monitor fifo_monitor_235;
    df_fifo_intf fifo_intf_236(clock,reset);
    assign fifo_intf_236.rd_en = AESL_inst_myproject.layer2_out_235_U.if_read & AESL_inst_myproject.layer2_out_235_U.if_empty_n;
    assign fifo_intf_236.wr_en = AESL_inst_myproject.layer2_out_235_U.if_write & AESL_inst_myproject.layer2_out_235_U.if_full_n;
    assign fifo_intf_236.fifo_rd_block = 0;
    assign fifo_intf_236.fifo_wr_block = 0;
    assign fifo_intf_236.finish = finish;
    csv_file_dump fifo_csv_dumper_236;
    csv_file_dump cstatus_csv_dumper_236;
    df_fifo_monitor fifo_monitor_236;
    df_fifo_intf fifo_intf_237(clock,reset);
    assign fifo_intf_237.rd_en = AESL_inst_myproject.layer2_out_236_U.if_read & AESL_inst_myproject.layer2_out_236_U.if_empty_n;
    assign fifo_intf_237.wr_en = AESL_inst_myproject.layer2_out_236_U.if_write & AESL_inst_myproject.layer2_out_236_U.if_full_n;
    assign fifo_intf_237.fifo_rd_block = 0;
    assign fifo_intf_237.fifo_wr_block = 0;
    assign fifo_intf_237.finish = finish;
    csv_file_dump fifo_csv_dumper_237;
    csv_file_dump cstatus_csv_dumper_237;
    df_fifo_monitor fifo_monitor_237;
    df_fifo_intf fifo_intf_238(clock,reset);
    assign fifo_intf_238.rd_en = AESL_inst_myproject.layer2_out_237_U.if_read & AESL_inst_myproject.layer2_out_237_U.if_empty_n;
    assign fifo_intf_238.wr_en = AESL_inst_myproject.layer2_out_237_U.if_write & AESL_inst_myproject.layer2_out_237_U.if_full_n;
    assign fifo_intf_238.fifo_rd_block = 0;
    assign fifo_intf_238.fifo_wr_block = 0;
    assign fifo_intf_238.finish = finish;
    csv_file_dump fifo_csv_dumper_238;
    csv_file_dump cstatus_csv_dumper_238;
    df_fifo_monitor fifo_monitor_238;
    df_fifo_intf fifo_intf_239(clock,reset);
    assign fifo_intf_239.rd_en = AESL_inst_myproject.layer2_out_238_U.if_read & AESL_inst_myproject.layer2_out_238_U.if_empty_n;
    assign fifo_intf_239.wr_en = AESL_inst_myproject.layer2_out_238_U.if_write & AESL_inst_myproject.layer2_out_238_U.if_full_n;
    assign fifo_intf_239.fifo_rd_block = 0;
    assign fifo_intf_239.fifo_wr_block = 0;
    assign fifo_intf_239.finish = finish;
    csv_file_dump fifo_csv_dumper_239;
    csv_file_dump cstatus_csv_dumper_239;
    df_fifo_monitor fifo_monitor_239;
    df_fifo_intf fifo_intf_240(clock,reset);
    assign fifo_intf_240.rd_en = AESL_inst_myproject.layer2_out_239_U.if_read & AESL_inst_myproject.layer2_out_239_U.if_empty_n;
    assign fifo_intf_240.wr_en = AESL_inst_myproject.layer2_out_239_U.if_write & AESL_inst_myproject.layer2_out_239_U.if_full_n;
    assign fifo_intf_240.fifo_rd_block = 0;
    assign fifo_intf_240.fifo_wr_block = 0;
    assign fifo_intf_240.finish = finish;
    csv_file_dump fifo_csv_dumper_240;
    csv_file_dump cstatus_csv_dumper_240;
    df_fifo_monitor fifo_monitor_240;
    df_fifo_intf fifo_intf_241(clock,reset);
    assign fifo_intf_241.rd_en = AESL_inst_myproject.layer2_out_240_U.if_read & AESL_inst_myproject.layer2_out_240_U.if_empty_n;
    assign fifo_intf_241.wr_en = AESL_inst_myproject.layer2_out_240_U.if_write & AESL_inst_myproject.layer2_out_240_U.if_full_n;
    assign fifo_intf_241.fifo_rd_block = 0;
    assign fifo_intf_241.fifo_wr_block = 0;
    assign fifo_intf_241.finish = finish;
    csv_file_dump fifo_csv_dumper_241;
    csv_file_dump cstatus_csv_dumper_241;
    df_fifo_monitor fifo_monitor_241;
    df_fifo_intf fifo_intf_242(clock,reset);
    assign fifo_intf_242.rd_en = AESL_inst_myproject.layer2_out_241_U.if_read & AESL_inst_myproject.layer2_out_241_U.if_empty_n;
    assign fifo_intf_242.wr_en = AESL_inst_myproject.layer2_out_241_U.if_write & AESL_inst_myproject.layer2_out_241_U.if_full_n;
    assign fifo_intf_242.fifo_rd_block = 0;
    assign fifo_intf_242.fifo_wr_block = 0;
    assign fifo_intf_242.finish = finish;
    csv_file_dump fifo_csv_dumper_242;
    csv_file_dump cstatus_csv_dumper_242;
    df_fifo_monitor fifo_monitor_242;
    df_fifo_intf fifo_intf_243(clock,reset);
    assign fifo_intf_243.rd_en = AESL_inst_myproject.layer2_out_242_U.if_read & AESL_inst_myproject.layer2_out_242_U.if_empty_n;
    assign fifo_intf_243.wr_en = AESL_inst_myproject.layer2_out_242_U.if_write & AESL_inst_myproject.layer2_out_242_U.if_full_n;
    assign fifo_intf_243.fifo_rd_block = 0;
    assign fifo_intf_243.fifo_wr_block = 0;
    assign fifo_intf_243.finish = finish;
    csv_file_dump fifo_csv_dumper_243;
    csv_file_dump cstatus_csv_dumper_243;
    df_fifo_monitor fifo_monitor_243;
    df_fifo_intf fifo_intf_244(clock,reset);
    assign fifo_intf_244.rd_en = AESL_inst_myproject.layer2_out_243_U.if_read & AESL_inst_myproject.layer2_out_243_U.if_empty_n;
    assign fifo_intf_244.wr_en = AESL_inst_myproject.layer2_out_243_U.if_write & AESL_inst_myproject.layer2_out_243_U.if_full_n;
    assign fifo_intf_244.fifo_rd_block = 0;
    assign fifo_intf_244.fifo_wr_block = 0;
    assign fifo_intf_244.finish = finish;
    csv_file_dump fifo_csv_dumper_244;
    csv_file_dump cstatus_csv_dumper_244;
    df_fifo_monitor fifo_monitor_244;
    df_fifo_intf fifo_intf_245(clock,reset);
    assign fifo_intf_245.rd_en = AESL_inst_myproject.layer2_out_244_U.if_read & AESL_inst_myproject.layer2_out_244_U.if_empty_n;
    assign fifo_intf_245.wr_en = AESL_inst_myproject.layer2_out_244_U.if_write & AESL_inst_myproject.layer2_out_244_U.if_full_n;
    assign fifo_intf_245.fifo_rd_block = 0;
    assign fifo_intf_245.fifo_wr_block = 0;
    assign fifo_intf_245.finish = finish;
    csv_file_dump fifo_csv_dumper_245;
    csv_file_dump cstatus_csv_dumper_245;
    df_fifo_monitor fifo_monitor_245;
    df_fifo_intf fifo_intf_246(clock,reset);
    assign fifo_intf_246.rd_en = AESL_inst_myproject.layer2_out_245_U.if_read & AESL_inst_myproject.layer2_out_245_U.if_empty_n;
    assign fifo_intf_246.wr_en = AESL_inst_myproject.layer2_out_245_U.if_write & AESL_inst_myproject.layer2_out_245_U.if_full_n;
    assign fifo_intf_246.fifo_rd_block = 0;
    assign fifo_intf_246.fifo_wr_block = 0;
    assign fifo_intf_246.finish = finish;
    csv_file_dump fifo_csv_dumper_246;
    csv_file_dump cstatus_csv_dumper_246;
    df_fifo_monitor fifo_monitor_246;
    df_fifo_intf fifo_intf_247(clock,reset);
    assign fifo_intf_247.rd_en = AESL_inst_myproject.layer2_out_246_U.if_read & AESL_inst_myproject.layer2_out_246_U.if_empty_n;
    assign fifo_intf_247.wr_en = AESL_inst_myproject.layer2_out_246_U.if_write & AESL_inst_myproject.layer2_out_246_U.if_full_n;
    assign fifo_intf_247.fifo_rd_block = 0;
    assign fifo_intf_247.fifo_wr_block = 0;
    assign fifo_intf_247.finish = finish;
    csv_file_dump fifo_csv_dumper_247;
    csv_file_dump cstatus_csv_dumper_247;
    df_fifo_monitor fifo_monitor_247;
    df_fifo_intf fifo_intf_248(clock,reset);
    assign fifo_intf_248.rd_en = AESL_inst_myproject.layer2_out_247_U.if_read & AESL_inst_myproject.layer2_out_247_U.if_empty_n;
    assign fifo_intf_248.wr_en = AESL_inst_myproject.layer2_out_247_U.if_write & AESL_inst_myproject.layer2_out_247_U.if_full_n;
    assign fifo_intf_248.fifo_rd_block = 0;
    assign fifo_intf_248.fifo_wr_block = 0;
    assign fifo_intf_248.finish = finish;
    csv_file_dump fifo_csv_dumper_248;
    csv_file_dump cstatus_csv_dumper_248;
    df_fifo_monitor fifo_monitor_248;
    df_fifo_intf fifo_intf_249(clock,reset);
    assign fifo_intf_249.rd_en = AESL_inst_myproject.layer2_out_248_U.if_read & AESL_inst_myproject.layer2_out_248_U.if_empty_n;
    assign fifo_intf_249.wr_en = AESL_inst_myproject.layer2_out_248_U.if_write & AESL_inst_myproject.layer2_out_248_U.if_full_n;
    assign fifo_intf_249.fifo_rd_block = 0;
    assign fifo_intf_249.fifo_wr_block = 0;
    assign fifo_intf_249.finish = finish;
    csv_file_dump fifo_csv_dumper_249;
    csv_file_dump cstatus_csv_dumper_249;
    df_fifo_monitor fifo_monitor_249;
    df_fifo_intf fifo_intf_250(clock,reset);
    assign fifo_intf_250.rd_en = AESL_inst_myproject.layer2_out_249_U.if_read & AESL_inst_myproject.layer2_out_249_U.if_empty_n;
    assign fifo_intf_250.wr_en = AESL_inst_myproject.layer2_out_249_U.if_write & AESL_inst_myproject.layer2_out_249_U.if_full_n;
    assign fifo_intf_250.fifo_rd_block = 0;
    assign fifo_intf_250.fifo_wr_block = 0;
    assign fifo_intf_250.finish = finish;
    csv_file_dump fifo_csv_dumper_250;
    csv_file_dump cstatus_csv_dumper_250;
    df_fifo_monitor fifo_monitor_250;
    df_fifo_intf fifo_intf_251(clock,reset);
    assign fifo_intf_251.rd_en = AESL_inst_myproject.layer2_out_250_U.if_read & AESL_inst_myproject.layer2_out_250_U.if_empty_n;
    assign fifo_intf_251.wr_en = AESL_inst_myproject.layer2_out_250_U.if_write & AESL_inst_myproject.layer2_out_250_U.if_full_n;
    assign fifo_intf_251.fifo_rd_block = 0;
    assign fifo_intf_251.fifo_wr_block = 0;
    assign fifo_intf_251.finish = finish;
    csv_file_dump fifo_csv_dumper_251;
    csv_file_dump cstatus_csv_dumper_251;
    df_fifo_monitor fifo_monitor_251;
    df_fifo_intf fifo_intf_252(clock,reset);
    assign fifo_intf_252.rd_en = AESL_inst_myproject.layer2_out_251_U.if_read & AESL_inst_myproject.layer2_out_251_U.if_empty_n;
    assign fifo_intf_252.wr_en = AESL_inst_myproject.layer2_out_251_U.if_write & AESL_inst_myproject.layer2_out_251_U.if_full_n;
    assign fifo_intf_252.fifo_rd_block = 0;
    assign fifo_intf_252.fifo_wr_block = 0;
    assign fifo_intf_252.finish = finish;
    csv_file_dump fifo_csv_dumper_252;
    csv_file_dump cstatus_csv_dumper_252;
    df_fifo_monitor fifo_monitor_252;
    df_fifo_intf fifo_intf_253(clock,reset);
    assign fifo_intf_253.rd_en = AESL_inst_myproject.layer2_out_252_U.if_read & AESL_inst_myproject.layer2_out_252_U.if_empty_n;
    assign fifo_intf_253.wr_en = AESL_inst_myproject.layer2_out_252_U.if_write & AESL_inst_myproject.layer2_out_252_U.if_full_n;
    assign fifo_intf_253.fifo_rd_block = 0;
    assign fifo_intf_253.fifo_wr_block = 0;
    assign fifo_intf_253.finish = finish;
    csv_file_dump fifo_csv_dumper_253;
    csv_file_dump cstatus_csv_dumper_253;
    df_fifo_monitor fifo_monitor_253;
    df_fifo_intf fifo_intf_254(clock,reset);
    assign fifo_intf_254.rd_en = AESL_inst_myproject.layer2_out_253_U.if_read & AESL_inst_myproject.layer2_out_253_U.if_empty_n;
    assign fifo_intf_254.wr_en = AESL_inst_myproject.layer2_out_253_U.if_write & AESL_inst_myproject.layer2_out_253_U.if_full_n;
    assign fifo_intf_254.fifo_rd_block = 0;
    assign fifo_intf_254.fifo_wr_block = 0;
    assign fifo_intf_254.finish = finish;
    csv_file_dump fifo_csv_dumper_254;
    csv_file_dump cstatus_csv_dumper_254;
    df_fifo_monitor fifo_monitor_254;
    df_fifo_intf fifo_intf_255(clock,reset);
    assign fifo_intf_255.rd_en = AESL_inst_myproject.layer2_out_254_U.if_read & AESL_inst_myproject.layer2_out_254_U.if_empty_n;
    assign fifo_intf_255.wr_en = AESL_inst_myproject.layer2_out_254_U.if_write & AESL_inst_myproject.layer2_out_254_U.if_full_n;
    assign fifo_intf_255.fifo_rd_block = 0;
    assign fifo_intf_255.fifo_wr_block = 0;
    assign fifo_intf_255.finish = finish;
    csv_file_dump fifo_csv_dumper_255;
    csv_file_dump cstatus_csv_dumper_255;
    df_fifo_monitor fifo_monitor_255;
    df_fifo_intf fifo_intf_256(clock,reset);
    assign fifo_intf_256.rd_en = AESL_inst_myproject.layer2_out_255_U.if_read & AESL_inst_myproject.layer2_out_255_U.if_empty_n;
    assign fifo_intf_256.wr_en = AESL_inst_myproject.layer2_out_255_U.if_write & AESL_inst_myproject.layer2_out_255_U.if_full_n;
    assign fifo_intf_256.fifo_rd_block = 0;
    assign fifo_intf_256.fifo_wr_block = 0;
    assign fifo_intf_256.finish = finish;
    csv_file_dump fifo_csv_dumper_256;
    csv_file_dump cstatus_csv_dumper_256;
    df_fifo_monitor fifo_monitor_256;
    df_fifo_intf fifo_intf_257(clock,reset);
    assign fifo_intf_257.rd_en = AESL_inst_myproject.layer2_out_256_U.if_read & AESL_inst_myproject.layer2_out_256_U.if_empty_n;
    assign fifo_intf_257.wr_en = AESL_inst_myproject.layer2_out_256_U.if_write & AESL_inst_myproject.layer2_out_256_U.if_full_n;
    assign fifo_intf_257.fifo_rd_block = 0;
    assign fifo_intf_257.fifo_wr_block = 0;
    assign fifo_intf_257.finish = finish;
    csv_file_dump fifo_csv_dumper_257;
    csv_file_dump cstatus_csv_dumper_257;
    df_fifo_monitor fifo_monitor_257;
    df_fifo_intf fifo_intf_258(clock,reset);
    assign fifo_intf_258.rd_en = AESL_inst_myproject.layer2_out_257_U.if_read & AESL_inst_myproject.layer2_out_257_U.if_empty_n;
    assign fifo_intf_258.wr_en = AESL_inst_myproject.layer2_out_257_U.if_write & AESL_inst_myproject.layer2_out_257_U.if_full_n;
    assign fifo_intf_258.fifo_rd_block = 0;
    assign fifo_intf_258.fifo_wr_block = 0;
    assign fifo_intf_258.finish = finish;
    csv_file_dump fifo_csv_dumper_258;
    csv_file_dump cstatus_csv_dumper_258;
    df_fifo_monitor fifo_monitor_258;
    df_fifo_intf fifo_intf_259(clock,reset);
    assign fifo_intf_259.rd_en = AESL_inst_myproject.layer2_out_258_U.if_read & AESL_inst_myproject.layer2_out_258_U.if_empty_n;
    assign fifo_intf_259.wr_en = AESL_inst_myproject.layer2_out_258_U.if_write & AESL_inst_myproject.layer2_out_258_U.if_full_n;
    assign fifo_intf_259.fifo_rd_block = 0;
    assign fifo_intf_259.fifo_wr_block = 0;
    assign fifo_intf_259.finish = finish;
    csv_file_dump fifo_csv_dumper_259;
    csv_file_dump cstatus_csv_dumper_259;
    df_fifo_monitor fifo_monitor_259;
    df_fifo_intf fifo_intf_260(clock,reset);
    assign fifo_intf_260.rd_en = AESL_inst_myproject.layer2_out_259_U.if_read & AESL_inst_myproject.layer2_out_259_U.if_empty_n;
    assign fifo_intf_260.wr_en = AESL_inst_myproject.layer2_out_259_U.if_write & AESL_inst_myproject.layer2_out_259_U.if_full_n;
    assign fifo_intf_260.fifo_rd_block = 0;
    assign fifo_intf_260.fifo_wr_block = 0;
    assign fifo_intf_260.finish = finish;
    csv_file_dump fifo_csv_dumper_260;
    csv_file_dump cstatus_csv_dumper_260;
    df_fifo_monitor fifo_monitor_260;
    df_fifo_intf fifo_intf_261(clock,reset);
    assign fifo_intf_261.rd_en = AESL_inst_myproject.layer2_out_260_U.if_read & AESL_inst_myproject.layer2_out_260_U.if_empty_n;
    assign fifo_intf_261.wr_en = AESL_inst_myproject.layer2_out_260_U.if_write & AESL_inst_myproject.layer2_out_260_U.if_full_n;
    assign fifo_intf_261.fifo_rd_block = 0;
    assign fifo_intf_261.fifo_wr_block = 0;
    assign fifo_intf_261.finish = finish;
    csv_file_dump fifo_csv_dumper_261;
    csv_file_dump cstatus_csv_dumper_261;
    df_fifo_monitor fifo_monitor_261;
    df_fifo_intf fifo_intf_262(clock,reset);
    assign fifo_intf_262.rd_en = AESL_inst_myproject.layer2_out_261_U.if_read & AESL_inst_myproject.layer2_out_261_U.if_empty_n;
    assign fifo_intf_262.wr_en = AESL_inst_myproject.layer2_out_261_U.if_write & AESL_inst_myproject.layer2_out_261_U.if_full_n;
    assign fifo_intf_262.fifo_rd_block = 0;
    assign fifo_intf_262.fifo_wr_block = 0;
    assign fifo_intf_262.finish = finish;
    csv_file_dump fifo_csv_dumper_262;
    csv_file_dump cstatus_csv_dumper_262;
    df_fifo_monitor fifo_monitor_262;
    df_fifo_intf fifo_intf_263(clock,reset);
    assign fifo_intf_263.rd_en = AESL_inst_myproject.layer2_out_262_U.if_read & AESL_inst_myproject.layer2_out_262_U.if_empty_n;
    assign fifo_intf_263.wr_en = AESL_inst_myproject.layer2_out_262_U.if_write & AESL_inst_myproject.layer2_out_262_U.if_full_n;
    assign fifo_intf_263.fifo_rd_block = 0;
    assign fifo_intf_263.fifo_wr_block = 0;
    assign fifo_intf_263.finish = finish;
    csv_file_dump fifo_csv_dumper_263;
    csv_file_dump cstatus_csv_dumper_263;
    df_fifo_monitor fifo_monitor_263;
    df_fifo_intf fifo_intf_264(clock,reset);
    assign fifo_intf_264.rd_en = AESL_inst_myproject.layer2_out_263_U.if_read & AESL_inst_myproject.layer2_out_263_U.if_empty_n;
    assign fifo_intf_264.wr_en = AESL_inst_myproject.layer2_out_263_U.if_write & AESL_inst_myproject.layer2_out_263_U.if_full_n;
    assign fifo_intf_264.fifo_rd_block = 0;
    assign fifo_intf_264.fifo_wr_block = 0;
    assign fifo_intf_264.finish = finish;
    csv_file_dump fifo_csv_dumper_264;
    csv_file_dump cstatus_csv_dumper_264;
    df_fifo_monitor fifo_monitor_264;
    df_fifo_intf fifo_intf_265(clock,reset);
    assign fifo_intf_265.rd_en = AESL_inst_myproject.layer2_out_264_U.if_read & AESL_inst_myproject.layer2_out_264_U.if_empty_n;
    assign fifo_intf_265.wr_en = AESL_inst_myproject.layer2_out_264_U.if_write & AESL_inst_myproject.layer2_out_264_U.if_full_n;
    assign fifo_intf_265.fifo_rd_block = 0;
    assign fifo_intf_265.fifo_wr_block = 0;
    assign fifo_intf_265.finish = finish;
    csv_file_dump fifo_csv_dumper_265;
    csv_file_dump cstatus_csv_dumper_265;
    df_fifo_monitor fifo_monitor_265;
    df_fifo_intf fifo_intf_266(clock,reset);
    assign fifo_intf_266.rd_en = AESL_inst_myproject.layer2_out_265_U.if_read & AESL_inst_myproject.layer2_out_265_U.if_empty_n;
    assign fifo_intf_266.wr_en = AESL_inst_myproject.layer2_out_265_U.if_write & AESL_inst_myproject.layer2_out_265_U.if_full_n;
    assign fifo_intf_266.fifo_rd_block = 0;
    assign fifo_intf_266.fifo_wr_block = 0;
    assign fifo_intf_266.finish = finish;
    csv_file_dump fifo_csv_dumper_266;
    csv_file_dump cstatus_csv_dumper_266;
    df_fifo_monitor fifo_monitor_266;
    df_fifo_intf fifo_intf_267(clock,reset);
    assign fifo_intf_267.rd_en = AESL_inst_myproject.layer2_out_266_U.if_read & AESL_inst_myproject.layer2_out_266_U.if_empty_n;
    assign fifo_intf_267.wr_en = AESL_inst_myproject.layer2_out_266_U.if_write & AESL_inst_myproject.layer2_out_266_U.if_full_n;
    assign fifo_intf_267.fifo_rd_block = 0;
    assign fifo_intf_267.fifo_wr_block = 0;
    assign fifo_intf_267.finish = finish;
    csv_file_dump fifo_csv_dumper_267;
    csv_file_dump cstatus_csv_dumper_267;
    df_fifo_monitor fifo_monitor_267;
    df_fifo_intf fifo_intf_268(clock,reset);
    assign fifo_intf_268.rd_en = AESL_inst_myproject.layer2_out_267_U.if_read & AESL_inst_myproject.layer2_out_267_U.if_empty_n;
    assign fifo_intf_268.wr_en = AESL_inst_myproject.layer2_out_267_U.if_write & AESL_inst_myproject.layer2_out_267_U.if_full_n;
    assign fifo_intf_268.fifo_rd_block = 0;
    assign fifo_intf_268.fifo_wr_block = 0;
    assign fifo_intf_268.finish = finish;
    csv_file_dump fifo_csv_dumper_268;
    csv_file_dump cstatus_csv_dumper_268;
    df_fifo_monitor fifo_monitor_268;
    df_fifo_intf fifo_intf_269(clock,reset);
    assign fifo_intf_269.rd_en = AESL_inst_myproject.layer2_out_268_U.if_read & AESL_inst_myproject.layer2_out_268_U.if_empty_n;
    assign fifo_intf_269.wr_en = AESL_inst_myproject.layer2_out_268_U.if_write & AESL_inst_myproject.layer2_out_268_U.if_full_n;
    assign fifo_intf_269.fifo_rd_block = 0;
    assign fifo_intf_269.fifo_wr_block = 0;
    assign fifo_intf_269.finish = finish;
    csv_file_dump fifo_csv_dumper_269;
    csv_file_dump cstatus_csv_dumper_269;
    df_fifo_monitor fifo_monitor_269;
    df_fifo_intf fifo_intf_270(clock,reset);
    assign fifo_intf_270.rd_en = AESL_inst_myproject.layer2_out_269_U.if_read & AESL_inst_myproject.layer2_out_269_U.if_empty_n;
    assign fifo_intf_270.wr_en = AESL_inst_myproject.layer2_out_269_U.if_write & AESL_inst_myproject.layer2_out_269_U.if_full_n;
    assign fifo_intf_270.fifo_rd_block = 0;
    assign fifo_intf_270.fifo_wr_block = 0;
    assign fifo_intf_270.finish = finish;
    csv_file_dump fifo_csv_dumper_270;
    csv_file_dump cstatus_csv_dumper_270;
    df_fifo_monitor fifo_monitor_270;
    df_fifo_intf fifo_intf_271(clock,reset);
    assign fifo_intf_271.rd_en = AESL_inst_myproject.layer2_out_270_U.if_read & AESL_inst_myproject.layer2_out_270_U.if_empty_n;
    assign fifo_intf_271.wr_en = AESL_inst_myproject.layer2_out_270_U.if_write & AESL_inst_myproject.layer2_out_270_U.if_full_n;
    assign fifo_intf_271.fifo_rd_block = 0;
    assign fifo_intf_271.fifo_wr_block = 0;
    assign fifo_intf_271.finish = finish;
    csv_file_dump fifo_csv_dumper_271;
    csv_file_dump cstatus_csv_dumper_271;
    df_fifo_monitor fifo_monitor_271;
    df_fifo_intf fifo_intf_272(clock,reset);
    assign fifo_intf_272.rd_en = AESL_inst_myproject.layer2_out_271_U.if_read & AESL_inst_myproject.layer2_out_271_U.if_empty_n;
    assign fifo_intf_272.wr_en = AESL_inst_myproject.layer2_out_271_U.if_write & AESL_inst_myproject.layer2_out_271_U.if_full_n;
    assign fifo_intf_272.fifo_rd_block = 0;
    assign fifo_intf_272.fifo_wr_block = 0;
    assign fifo_intf_272.finish = finish;
    csv_file_dump fifo_csv_dumper_272;
    csv_file_dump cstatus_csv_dumper_272;
    df_fifo_monitor fifo_monitor_272;
    df_fifo_intf fifo_intf_273(clock,reset);
    assign fifo_intf_273.rd_en = AESL_inst_myproject.layer2_out_272_U.if_read & AESL_inst_myproject.layer2_out_272_U.if_empty_n;
    assign fifo_intf_273.wr_en = AESL_inst_myproject.layer2_out_272_U.if_write & AESL_inst_myproject.layer2_out_272_U.if_full_n;
    assign fifo_intf_273.fifo_rd_block = 0;
    assign fifo_intf_273.fifo_wr_block = 0;
    assign fifo_intf_273.finish = finish;
    csv_file_dump fifo_csv_dumper_273;
    csv_file_dump cstatus_csv_dumper_273;
    df_fifo_monitor fifo_monitor_273;
    df_fifo_intf fifo_intf_274(clock,reset);
    assign fifo_intf_274.rd_en = AESL_inst_myproject.layer2_out_273_U.if_read & AESL_inst_myproject.layer2_out_273_U.if_empty_n;
    assign fifo_intf_274.wr_en = AESL_inst_myproject.layer2_out_273_U.if_write & AESL_inst_myproject.layer2_out_273_U.if_full_n;
    assign fifo_intf_274.fifo_rd_block = 0;
    assign fifo_intf_274.fifo_wr_block = 0;
    assign fifo_intf_274.finish = finish;
    csv_file_dump fifo_csv_dumper_274;
    csv_file_dump cstatus_csv_dumper_274;
    df_fifo_monitor fifo_monitor_274;
    df_fifo_intf fifo_intf_275(clock,reset);
    assign fifo_intf_275.rd_en = AESL_inst_myproject.layer2_out_274_U.if_read & AESL_inst_myproject.layer2_out_274_U.if_empty_n;
    assign fifo_intf_275.wr_en = AESL_inst_myproject.layer2_out_274_U.if_write & AESL_inst_myproject.layer2_out_274_U.if_full_n;
    assign fifo_intf_275.fifo_rd_block = 0;
    assign fifo_intf_275.fifo_wr_block = 0;
    assign fifo_intf_275.finish = finish;
    csv_file_dump fifo_csv_dumper_275;
    csv_file_dump cstatus_csv_dumper_275;
    df_fifo_monitor fifo_monitor_275;
    df_fifo_intf fifo_intf_276(clock,reset);
    assign fifo_intf_276.rd_en = AESL_inst_myproject.layer2_out_275_U.if_read & AESL_inst_myproject.layer2_out_275_U.if_empty_n;
    assign fifo_intf_276.wr_en = AESL_inst_myproject.layer2_out_275_U.if_write & AESL_inst_myproject.layer2_out_275_U.if_full_n;
    assign fifo_intf_276.fifo_rd_block = 0;
    assign fifo_intf_276.fifo_wr_block = 0;
    assign fifo_intf_276.finish = finish;
    csv_file_dump fifo_csv_dumper_276;
    csv_file_dump cstatus_csv_dumper_276;
    df_fifo_monitor fifo_monitor_276;
    df_fifo_intf fifo_intf_277(clock,reset);
    assign fifo_intf_277.rd_en = AESL_inst_myproject.layer2_out_276_U.if_read & AESL_inst_myproject.layer2_out_276_U.if_empty_n;
    assign fifo_intf_277.wr_en = AESL_inst_myproject.layer2_out_276_U.if_write & AESL_inst_myproject.layer2_out_276_U.if_full_n;
    assign fifo_intf_277.fifo_rd_block = 0;
    assign fifo_intf_277.fifo_wr_block = 0;
    assign fifo_intf_277.finish = finish;
    csv_file_dump fifo_csv_dumper_277;
    csv_file_dump cstatus_csv_dumper_277;
    df_fifo_monitor fifo_monitor_277;
    df_fifo_intf fifo_intf_278(clock,reset);
    assign fifo_intf_278.rd_en = AESL_inst_myproject.layer2_out_277_U.if_read & AESL_inst_myproject.layer2_out_277_U.if_empty_n;
    assign fifo_intf_278.wr_en = AESL_inst_myproject.layer2_out_277_U.if_write & AESL_inst_myproject.layer2_out_277_U.if_full_n;
    assign fifo_intf_278.fifo_rd_block = 0;
    assign fifo_intf_278.fifo_wr_block = 0;
    assign fifo_intf_278.finish = finish;
    csv_file_dump fifo_csv_dumper_278;
    csv_file_dump cstatus_csv_dumper_278;
    df_fifo_monitor fifo_monitor_278;
    df_fifo_intf fifo_intf_279(clock,reset);
    assign fifo_intf_279.rd_en = AESL_inst_myproject.layer2_out_278_U.if_read & AESL_inst_myproject.layer2_out_278_U.if_empty_n;
    assign fifo_intf_279.wr_en = AESL_inst_myproject.layer2_out_278_U.if_write & AESL_inst_myproject.layer2_out_278_U.if_full_n;
    assign fifo_intf_279.fifo_rd_block = 0;
    assign fifo_intf_279.fifo_wr_block = 0;
    assign fifo_intf_279.finish = finish;
    csv_file_dump fifo_csv_dumper_279;
    csv_file_dump cstatus_csv_dumper_279;
    df_fifo_monitor fifo_monitor_279;
    df_fifo_intf fifo_intf_280(clock,reset);
    assign fifo_intf_280.rd_en = AESL_inst_myproject.layer2_out_279_U.if_read & AESL_inst_myproject.layer2_out_279_U.if_empty_n;
    assign fifo_intf_280.wr_en = AESL_inst_myproject.layer2_out_279_U.if_write & AESL_inst_myproject.layer2_out_279_U.if_full_n;
    assign fifo_intf_280.fifo_rd_block = 0;
    assign fifo_intf_280.fifo_wr_block = 0;
    assign fifo_intf_280.finish = finish;
    csv_file_dump fifo_csv_dumper_280;
    csv_file_dump cstatus_csv_dumper_280;
    df_fifo_monitor fifo_monitor_280;
    df_fifo_intf fifo_intf_281(clock,reset);
    assign fifo_intf_281.rd_en = AESL_inst_myproject.layer2_out_280_U.if_read & AESL_inst_myproject.layer2_out_280_U.if_empty_n;
    assign fifo_intf_281.wr_en = AESL_inst_myproject.layer2_out_280_U.if_write & AESL_inst_myproject.layer2_out_280_U.if_full_n;
    assign fifo_intf_281.fifo_rd_block = 0;
    assign fifo_intf_281.fifo_wr_block = 0;
    assign fifo_intf_281.finish = finish;
    csv_file_dump fifo_csv_dumper_281;
    csv_file_dump cstatus_csv_dumper_281;
    df_fifo_monitor fifo_monitor_281;
    df_fifo_intf fifo_intf_282(clock,reset);
    assign fifo_intf_282.rd_en = AESL_inst_myproject.layer2_out_281_U.if_read & AESL_inst_myproject.layer2_out_281_U.if_empty_n;
    assign fifo_intf_282.wr_en = AESL_inst_myproject.layer2_out_281_U.if_write & AESL_inst_myproject.layer2_out_281_U.if_full_n;
    assign fifo_intf_282.fifo_rd_block = 0;
    assign fifo_intf_282.fifo_wr_block = 0;
    assign fifo_intf_282.finish = finish;
    csv_file_dump fifo_csv_dumper_282;
    csv_file_dump cstatus_csv_dumper_282;
    df_fifo_monitor fifo_monitor_282;
    df_fifo_intf fifo_intf_283(clock,reset);
    assign fifo_intf_283.rd_en = AESL_inst_myproject.layer2_out_282_U.if_read & AESL_inst_myproject.layer2_out_282_U.if_empty_n;
    assign fifo_intf_283.wr_en = AESL_inst_myproject.layer2_out_282_U.if_write & AESL_inst_myproject.layer2_out_282_U.if_full_n;
    assign fifo_intf_283.fifo_rd_block = 0;
    assign fifo_intf_283.fifo_wr_block = 0;
    assign fifo_intf_283.finish = finish;
    csv_file_dump fifo_csv_dumper_283;
    csv_file_dump cstatus_csv_dumper_283;
    df_fifo_monitor fifo_monitor_283;
    df_fifo_intf fifo_intf_284(clock,reset);
    assign fifo_intf_284.rd_en = AESL_inst_myproject.layer2_out_283_U.if_read & AESL_inst_myproject.layer2_out_283_U.if_empty_n;
    assign fifo_intf_284.wr_en = AESL_inst_myproject.layer2_out_283_U.if_write & AESL_inst_myproject.layer2_out_283_U.if_full_n;
    assign fifo_intf_284.fifo_rd_block = 0;
    assign fifo_intf_284.fifo_wr_block = 0;
    assign fifo_intf_284.finish = finish;
    csv_file_dump fifo_csv_dumper_284;
    csv_file_dump cstatus_csv_dumper_284;
    df_fifo_monitor fifo_monitor_284;
    df_fifo_intf fifo_intf_285(clock,reset);
    assign fifo_intf_285.rd_en = AESL_inst_myproject.layer2_out_284_U.if_read & AESL_inst_myproject.layer2_out_284_U.if_empty_n;
    assign fifo_intf_285.wr_en = AESL_inst_myproject.layer2_out_284_U.if_write & AESL_inst_myproject.layer2_out_284_U.if_full_n;
    assign fifo_intf_285.fifo_rd_block = 0;
    assign fifo_intf_285.fifo_wr_block = 0;
    assign fifo_intf_285.finish = finish;
    csv_file_dump fifo_csv_dumper_285;
    csv_file_dump cstatus_csv_dumper_285;
    df_fifo_monitor fifo_monitor_285;
    df_fifo_intf fifo_intf_286(clock,reset);
    assign fifo_intf_286.rd_en = AESL_inst_myproject.layer2_out_285_U.if_read & AESL_inst_myproject.layer2_out_285_U.if_empty_n;
    assign fifo_intf_286.wr_en = AESL_inst_myproject.layer2_out_285_U.if_write & AESL_inst_myproject.layer2_out_285_U.if_full_n;
    assign fifo_intf_286.fifo_rd_block = 0;
    assign fifo_intf_286.fifo_wr_block = 0;
    assign fifo_intf_286.finish = finish;
    csv_file_dump fifo_csv_dumper_286;
    csv_file_dump cstatus_csv_dumper_286;
    df_fifo_monitor fifo_monitor_286;
    df_fifo_intf fifo_intf_287(clock,reset);
    assign fifo_intf_287.rd_en = AESL_inst_myproject.layer2_out_286_U.if_read & AESL_inst_myproject.layer2_out_286_U.if_empty_n;
    assign fifo_intf_287.wr_en = AESL_inst_myproject.layer2_out_286_U.if_write & AESL_inst_myproject.layer2_out_286_U.if_full_n;
    assign fifo_intf_287.fifo_rd_block = 0;
    assign fifo_intf_287.fifo_wr_block = 0;
    assign fifo_intf_287.finish = finish;
    csv_file_dump fifo_csv_dumper_287;
    csv_file_dump cstatus_csv_dumper_287;
    df_fifo_monitor fifo_monitor_287;
    df_fifo_intf fifo_intf_288(clock,reset);
    assign fifo_intf_288.rd_en = AESL_inst_myproject.layer2_out_287_U.if_read & AESL_inst_myproject.layer2_out_287_U.if_empty_n;
    assign fifo_intf_288.wr_en = AESL_inst_myproject.layer2_out_287_U.if_write & AESL_inst_myproject.layer2_out_287_U.if_full_n;
    assign fifo_intf_288.fifo_rd_block = 0;
    assign fifo_intf_288.fifo_wr_block = 0;
    assign fifo_intf_288.finish = finish;
    csv_file_dump fifo_csv_dumper_288;
    csv_file_dump cstatus_csv_dumper_288;
    df_fifo_monitor fifo_monitor_288;
    df_fifo_intf fifo_intf_289(clock,reset);
    assign fifo_intf_289.rd_en = AESL_inst_myproject.layer2_out_288_U.if_read & AESL_inst_myproject.layer2_out_288_U.if_empty_n;
    assign fifo_intf_289.wr_en = AESL_inst_myproject.layer2_out_288_U.if_write & AESL_inst_myproject.layer2_out_288_U.if_full_n;
    assign fifo_intf_289.fifo_rd_block = 0;
    assign fifo_intf_289.fifo_wr_block = 0;
    assign fifo_intf_289.finish = finish;
    csv_file_dump fifo_csv_dumper_289;
    csv_file_dump cstatus_csv_dumper_289;
    df_fifo_monitor fifo_monitor_289;
    df_fifo_intf fifo_intf_290(clock,reset);
    assign fifo_intf_290.rd_en = AESL_inst_myproject.layer2_out_289_U.if_read & AESL_inst_myproject.layer2_out_289_U.if_empty_n;
    assign fifo_intf_290.wr_en = AESL_inst_myproject.layer2_out_289_U.if_write & AESL_inst_myproject.layer2_out_289_U.if_full_n;
    assign fifo_intf_290.fifo_rd_block = 0;
    assign fifo_intf_290.fifo_wr_block = 0;
    assign fifo_intf_290.finish = finish;
    csv_file_dump fifo_csv_dumper_290;
    csv_file_dump cstatus_csv_dumper_290;
    df_fifo_monitor fifo_monitor_290;
    df_fifo_intf fifo_intf_291(clock,reset);
    assign fifo_intf_291.rd_en = AESL_inst_myproject.layer2_out_290_U.if_read & AESL_inst_myproject.layer2_out_290_U.if_empty_n;
    assign fifo_intf_291.wr_en = AESL_inst_myproject.layer2_out_290_U.if_write & AESL_inst_myproject.layer2_out_290_U.if_full_n;
    assign fifo_intf_291.fifo_rd_block = 0;
    assign fifo_intf_291.fifo_wr_block = 0;
    assign fifo_intf_291.finish = finish;
    csv_file_dump fifo_csv_dumper_291;
    csv_file_dump cstatus_csv_dumper_291;
    df_fifo_monitor fifo_monitor_291;
    df_fifo_intf fifo_intf_292(clock,reset);
    assign fifo_intf_292.rd_en = AESL_inst_myproject.layer2_out_291_U.if_read & AESL_inst_myproject.layer2_out_291_U.if_empty_n;
    assign fifo_intf_292.wr_en = AESL_inst_myproject.layer2_out_291_U.if_write & AESL_inst_myproject.layer2_out_291_U.if_full_n;
    assign fifo_intf_292.fifo_rd_block = 0;
    assign fifo_intf_292.fifo_wr_block = 0;
    assign fifo_intf_292.finish = finish;
    csv_file_dump fifo_csv_dumper_292;
    csv_file_dump cstatus_csv_dumper_292;
    df_fifo_monitor fifo_monitor_292;
    df_fifo_intf fifo_intf_293(clock,reset);
    assign fifo_intf_293.rd_en = AESL_inst_myproject.layer2_out_292_U.if_read & AESL_inst_myproject.layer2_out_292_U.if_empty_n;
    assign fifo_intf_293.wr_en = AESL_inst_myproject.layer2_out_292_U.if_write & AESL_inst_myproject.layer2_out_292_U.if_full_n;
    assign fifo_intf_293.fifo_rd_block = 0;
    assign fifo_intf_293.fifo_wr_block = 0;
    assign fifo_intf_293.finish = finish;
    csv_file_dump fifo_csv_dumper_293;
    csv_file_dump cstatus_csv_dumper_293;
    df_fifo_monitor fifo_monitor_293;
    df_fifo_intf fifo_intf_294(clock,reset);
    assign fifo_intf_294.rd_en = AESL_inst_myproject.layer2_out_293_U.if_read & AESL_inst_myproject.layer2_out_293_U.if_empty_n;
    assign fifo_intf_294.wr_en = AESL_inst_myproject.layer2_out_293_U.if_write & AESL_inst_myproject.layer2_out_293_U.if_full_n;
    assign fifo_intf_294.fifo_rd_block = 0;
    assign fifo_intf_294.fifo_wr_block = 0;
    assign fifo_intf_294.finish = finish;
    csv_file_dump fifo_csv_dumper_294;
    csv_file_dump cstatus_csv_dumper_294;
    df_fifo_monitor fifo_monitor_294;
    df_fifo_intf fifo_intf_295(clock,reset);
    assign fifo_intf_295.rd_en = AESL_inst_myproject.layer2_out_294_U.if_read & AESL_inst_myproject.layer2_out_294_U.if_empty_n;
    assign fifo_intf_295.wr_en = AESL_inst_myproject.layer2_out_294_U.if_write & AESL_inst_myproject.layer2_out_294_U.if_full_n;
    assign fifo_intf_295.fifo_rd_block = 0;
    assign fifo_intf_295.fifo_wr_block = 0;
    assign fifo_intf_295.finish = finish;
    csv_file_dump fifo_csv_dumper_295;
    csv_file_dump cstatus_csv_dumper_295;
    df_fifo_monitor fifo_monitor_295;
    df_fifo_intf fifo_intf_296(clock,reset);
    assign fifo_intf_296.rd_en = AESL_inst_myproject.layer2_out_295_U.if_read & AESL_inst_myproject.layer2_out_295_U.if_empty_n;
    assign fifo_intf_296.wr_en = AESL_inst_myproject.layer2_out_295_U.if_write & AESL_inst_myproject.layer2_out_295_U.if_full_n;
    assign fifo_intf_296.fifo_rd_block = 0;
    assign fifo_intf_296.fifo_wr_block = 0;
    assign fifo_intf_296.finish = finish;
    csv_file_dump fifo_csv_dumper_296;
    csv_file_dump cstatus_csv_dumper_296;
    df_fifo_monitor fifo_monitor_296;
    df_fifo_intf fifo_intf_297(clock,reset);
    assign fifo_intf_297.rd_en = AESL_inst_myproject.layer2_out_296_U.if_read & AESL_inst_myproject.layer2_out_296_U.if_empty_n;
    assign fifo_intf_297.wr_en = AESL_inst_myproject.layer2_out_296_U.if_write & AESL_inst_myproject.layer2_out_296_U.if_full_n;
    assign fifo_intf_297.fifo_rd_block = 0;
    assign fifo_intf_297.fifo_wr_block = 0;
    assign fifo_intf_297.finish = finish;
    csv_file_dump fifo_csv_dumper_297;
    csv_file_dump cstatus_csv_dumper_297;
    df_fifo_monitor fifo_monitor_297;
    df_fifo_intf fifo_intf_298(clock,reset);
    assign fifo_intf_298.rd_en = AESL_inst_myproject.layer2_out_297_U.if_read & AESL_inst_myproject.layer2_out_297_U.if_empty_n;
    assign fifo_intf_298.wr_en = AESL_inst_myproject.layer2_out_297_U.if_write & AESL_inst_myproject.layer2_out_297_U.if_full_n;
    assign fifo_intf_298.fifo_rd_block = 0;
    assign fifo_intf_298.fifo_wr_block = 0;
    assign fifo_intf_298.finish = finish;
    csv_file_dump fifo_csv_dumper_298;
    csv_file_dump cstatus_csv_dumper_298;
    df_fifo_monitor fifo_monitor_298;
    df_fifo_intf fifo_intf_299(clock,reset);
    assign fifo_intf_299.rd_en = AESL_inst_myproject.layer2_out_298_U.if_read & AESL_inst_myproject.layer2_out_298_U.if_empty_n;
    assign fifo_intf_299.wr_en = AESL_inst_myproject.layer2_out_298_U.if_write & AESL_inst_myproject.layer2_out_298_U.if_full_n;
    assign fifo_intf_299.fifo_rd_block = 0;
    assign fifo_intf_299.fifo_wr_block = 0;
    assign fifo_intf_299.finish = finish;
    csv_file_dump fifo_csv_dumper_299;
    csv_file_dump cstatus_csv_dumper_299;
    df_fifo_monitor fifo_monitor_299;
    df_fifo_intf fifo_intf_300(clock,reset);
    assign fifo_intf_300.rd_en = AESL_inst_myproject.layer2_out_299_U.if_read & AESL_inst_myproject.layer2_out_299_U.if_empty_n;
    assign fifo_intf_300.wr_en = AESL_inst_myproject.layer2_out_299_U.if_write & AESL_inst_myproject.layer2_out_299_U.if_full_n;
    assign fifo_intf_300.fifo_rd_block = 0;
    assign fifo_intf_300.fifo_wr_block = 0;
    assign fifo_intf_300.finish = finish;
    csv_file_dump fifo_csv_dumper_300;
    csv_file_dump cstatus_csv_dumper_300;
    df_fifo_monitor fifo_monitor_300;
    df_fifo_intf fifo_intf_301(clock,reset);
    assign fifo_intf_301.rd_en = AESL_inst_myproject.layer2_out_300_U.if_read & AESL_inst_myproject.layer2_out_300_U.if_empty_n;
    assign fifo_intf_301.wr_en = AESL_inst_myproject.layer2_out_300_U.if_write & AESL_inst_myproject.layer2_out_300_U.if_full_n;
    assign fifo_intf_301.fifo_rd_block = 0;
    assign fifo_intf_301.fifo_wr_block = 0;
    assign fifo_intf_301.finish = finish;
    csv_file_dump fifo_csv_dumper_301;
    csv_file_dump cstatus_csv_dumper_301;
    df_fifo_monitor fifo_monitor_301;
    df_fifo_intf fifo_intf_302(clock,reset);
    assign fifo_intf_302.rd_en = AESL_inst_myproject.layer2_out_301_U.if_read & AESL_inst_myproject.layer2_out_301_U.if_empty_n;
    assign fifo_intf_302.wr_en = AESL_inst_myproject.layer2_out_301_U.if_write & AESL_inst_myproject.layer2_out_301_U.if_full_n;
    assign fifo_intf_302.fifo_rd_block = 0;
    assign fifo_intf_302.fifo_wr_block = 0;
    assign fifo_intf_302.finish = finish;
    csv_file_dump fifo_csv_dumper_302;
    csv_file_dump cstatus_csv_dumper_302;
    df_fifo_monitor fifo_monitor_302;
    df_fifo_intf fifo_intf_303(clock,reset);
    assign fifo_intf_303.rd_en = AESL_inst_myproject.layer2_out_302_U.if_read & AESL_inst_myproject.layer2_out_302_U.if_empty_n;
    assign fifo_intf_303.wr_en = AESL_inst_myproject.layer2_out_302_U.if_write & AESL_inst_myproject.layer2_out_302_U.if_full_n;
    assign fifo_intf_303.fifo_rd_block = 0;
    assign fifo_intf_303.fifo_wr_block = 0;
    assign fifo_intf_303.finish = finish;
    csv_file_dump fifo_csv_dumper_303;
    csv_file_dump cstatus_csv_dumper_303;
    df_fifo_monitor fifo_monitor_303;
    df_fifo_intf fifo_intf_304(clock,reset);
    assign fifo_intf_304.rd_en = AESL_inst_myproject.layer2_out_303_U.if_read & AESL_inst_myproject.layer2_out_303_U.if_empty_n;
    assign fifo_intf_304.wr_en = AESL_inst_myproject.layer2_out_303_U.if_write & AESL_inst_myproject.layer2_out_303_U.if_full_n;
    assign fifo_intf_304.fifo_rd_block = 0;
    assign fifo_intf_304.fifo_wr_block = 0;
    assign fifo_intf_304.finish = finish;
    csv_file_dump fifo_csv_dumper_304;
    csv_file_dump cstatus_csv_dumper_304;
    df_fifo_monitor fifo_monitor_304;
    df_fifo_intf fifo_intf_305(clock,reset);
    assign fifo_intf_305.rd_en = AESL_inst_myproject.layer2_out_304_U.if_read & AESL_inst_myproject.layer2_out_304_U.if_empty_n;
    assign fifo_intf_305.wr_en = AESL_inst_myproject.layer2_out_304_U.if_write & AESL_inst_myproject.layer2_out_304_U.if_full_n;
    assign fifo_intf_305.fifo_rd_block = 0;
    assign fifo_intf_305.fifo_wr_block = 0;
    assign fifo_intf_305.finish = finish;
    csv_file_dump fifo_csv_dumper_305;
    csv_file_dump cstatus_csv_dumper_305;
    df_fifo_monitor fifo_monitor_305;
    df_fifo_intf fifo_intf_306(clock,reset);
    assign fifo_intf_306.rd_en = AESL_inst_myproject.layer2_out_305_U.if_read & AESL_inst_myproject.layer2_out_305_U.if_empty_n;
    assign fifo_intf_306.wr_en = AESL_inst_myproject.layer2_out_305_U.if_write & AESL_inst_myproject.layer2_out_305_U.if_full_n;
    assign fifo_intf_306.fifo_rd_block = 0;
    assign fifo_intf_306.fifo_wr_block = 0;
    assign fifo_intf_306.finish = finish;
    csv_file_dump fifo_csv_dumper_306;
    csv_file_dump cstatus_csv_dumper_306;
    df_fifo_monitor fifo_monitor_306;
    df_fifo_intf fifo_intf_307(clock,reset);
    assign fifo_intf_307.rd_en = AESL_inst_myproject.layer2_out_306_U.if_read & AESL_inst_myproject.layer2_out_306_U.if_empty_n;
    assign fifo_intf_307.wr_en = AESL_inst_myproject.layer2_out_306_U.if_write & AESL_inst_myproject.layer2_out_306_U.if_full_n;
    assign fifo_intf_307.fifo_rd_block = 0;
    assign fifo_intf_307.fifo_wr_block = 0;
    assign fifo_intf_307.finish = finish;
    csv_file_dump fifo_csv_dumper_307;
    csv_file_dump cstatus_csv_dumper_307;
    df_fifo_monitor fifo_monitor_307;
    df_fifo_intf fifo_intf_308(clock,reset);
    assign fifo_intf_308.rd_en = AESL_inst_myproject.layer2_out_307_U.if_read & AESL_inst_myproject.layer2_out_307_U.if_empty_n;
    assign fifo_intf_308.wr_en = AESL_inst_myproject.layer2_out_307_U.if_write & AESL_inst_myproject.layer2_out_307_U.if_full_n;
    assign fifo_intf_308.fifo_rd_block = 0;
    assign fifo_intf_308.fifo_wr_block = 0;
    assign fifo_intf_308.finish = finish;
    csv_file_dump fifo_csv_dumper_308;
    csv_file_dump cstatus_csv_dumper_308;
    df_fifo_monitor fifo_monitor_308;
    df_fifo_intf fifo_intf_309(clock,reset);
    assign fifo_intf_309.rd_en = AESL_inst_myproject.layer2_out_308_U.if_read & AESL_inst_myproject.layer2_out_308_U.if_empty_n;
    assign fifo_intf_309.wr_en = AESL_inst_myproject.layer2_out_308_U.if_write & AESL_inst_myproject.layer2_out_308_U.if_full_n;
    assign fifo_intf_309.fifo_rd_block = 0;
    assign fifo_intf_309.fifo_wr_block = 0;
    assign fifo_intf_309.finish = finish;
    csv_file_dump fifo_csv_dumper_309;
    csv_file_dump cstatus_csv_dumper_309;
    df_fifo_monitor fifo_monitor_309;
    df_fifo_intf fifo_intf_310(clock,reset);
    assign fifo_intf_310.rd_en = AESL_inst_myproject.layer2_out_309_U.if_read & AESL_inst_myproject.layer2_out_309_U.if_empty_n;
    assign fifo_intf_310.wr_en = AESL_inst_myproject.layer2_out_309_U.if_write & AESL_inst_myproject.layer2_out_309_U.if_full_n;
    assign fifo_intf_310.fifo_rd_block = 0;
    assign fifo_intf_310.fifo_wr_block = 0;
    assign fifo_intf_310.finish = finish;
    csv_file_dump fifo_csv_dumper_310;
    csv_file_dump cstatus_csv_dumper_310;
    df_fifo_monitor fifo_monitor_310;
    df_fifo_intf fifo_intf_311(clock,reset);
    assign fifo_intf_311.rd_en = AESL_inst_myproject.layer2_out_310_U.if_read & AESL_inst_myproject.layer2_out_310_U.if_empty_n;
    assign fifo_intf_311.wr_en = AESL_inst_myproject.layer2_out_310_U.if_write & AESL_inst_myproject.layer2_out_310_U.if_full_n;
    assign fifo_intf_311.fifo_rd_block = 0;
    assign fifo_intf_311.fifo_wr_block = 0;
    assign fifo_intf_311.finish = finish;
    csv_file_dump fifo_csv_dumper_311;
    csv_file_dump cstatus_csv_dumper_311;
    df_fifo_monitor fifo_monitor_311;
    df_fifo_intf fifo_intf_312(clock,reset);
    assign fifo_intf_312.rd_en = AESL_inst_myproject.layer2_out_311_U.if_read & AESL_inst_myproject.layer2_out_311_U.if_empty_n;
    assign fifo_intf_312.wr_en = AESL_inst_myproject.layer2_out_311_U.if_write & AESL_inst_myproject.layer2_out_311_U.if_full_n;
    assign fifo_intf_312.fifo_rd_block = 0;
    assign fifo_intf_312.fifo_wr_block = 0;
    assign fifo_intf_312.finish = finish;
    csv_file_dump fifo_csv_dumper_312;
    csv_file_dump cstatus_csv_dumper_312;
    df_fifo_monitor fifo_monitor_312;
    df_fifo_intf fifo_intf_313(clock,reset);
    assign fifo_intf_313.rd_en = AESL_inst_myproject.layer2_out_312_U.if_read & AESL_inst_myproject.layer2_out_312_U.if_empty_n;
    assign fifo_intf_313.wr_en = AESL_inst_myproject.layer2_out_312_U.if_write & AESL_inst_myproject.layer2_out_312_U.if_full_n;
    assign fifo_intf_313.fifo_rd_block = 0;
    assign fifo_intf_313.fifo_wr_block = 0;
    assign fifo_intf_313.finish = finish;
    csv_file_dump fifo_csv_dumper_313;
    csv_file_dump cstatus_csv_dumper_313;
    df_fifo_monitor fifo_monitor_313;
    df_fifo_intf fifo_intf_314(clock,reset);
    assign fifo_intf_314.rd_en = AESL_inst_myproject.layer2_out_313_U.if_read & AESL_inst_myproject.layer2_out_313_U.if_empty_n;
    assign fifo_intf_314.wr_en = AESL_inst_myproject.layer2_out_313_U.if_write & AESL_inst_myproject.layer2_out_313_U.if_full_n;
    assign fifo_intf_314.fifo_rd_block = 0;
    assign fifo_intf_314.fifo_wr_block = 0;
    assign fifo_intf_314.finish = finish;
    csv_file_dump fifo_csv_dumper_314;
    csv_file_dump cstatus_csv_dumper_314;
    df_fifo_monitor fifo_monitor_314;
    df_fifo_intf fifo_intf_315(clock,reset);
    assign fifo_intf_315.rd_en = AESL_inst_myproject.layer2_out_314_U.if_read & AESL_inst_myproject.layer2_out_314_U.if_empty_n;
    assign fifo_intf_315.wr_en = AESL_inst_myproject.layer2_out_314_U.if_write & AESL_inst_myproject.layer2_out_314_U.if_full_n;
    assign fifo_intf_315.fifo_rd_block = 0;
    assign fifo_intf_315.fifo_wr_block = 0;
    assign fifo_intf_315.finish = finish;
    csv_file_dump fifo_csv_dumper_315;
    csv_file_dump cstatus_csv_dumper_315;
    df_fifo_monitor fifo_monitor_315;
    df_fifo_intf fifo_intf_316(clock,reset);
    assign fifo_intf_316.rd_en = AESL_inst_myproject.layer2_out_315_U.if_read & AESL_inst_myproject.layer2_out_315_U.if_empty_n;
    assign fifo_intf_316.wr_en = AESL_inst_myproject.layer2_out_315_U.if_write & AESL_inst_myproject.layer2_out_315_U.if_full_n;
    assign fifo_intf_316.fifo_rd_block = 0;
    assign fifo_intf_316.fifo_wr_block = 0;
    assign fifo_intf_316.finish = finish;
    csv_file_dump fifo_csv_dumper_316;
    csv_file_dump cstatus_csv_dumper_316;
    df_fifo_monitor fifo_monitor_316;
    df_fifo_intf fifo_intf_317(clock,reset);
    assign fifo_intf_317.rd_en = AESL_inst_myproject.layer2_out_316_U.if_read & AESL_inst_myproject.layer2_out_316_U.if_empty_n;
    assign fifo_intf_317.wr_en = AESL_inst_myproject.layer2_out_316_U.if_write & AESL_inst_myproject.layer2_out_316_U.if_full_n;
    assign fifo_intf_317.fifo_rd_block = 0;
    assign fifo_intf_317.fifo_wr_block = 0;
    assign fifo_intf_317.finish = finish;
    csv_file_dump fifo_csv_dumper_317;
    csv_file_dump cstatus_csv_dumper_317;
    df_fifo_monitor fifo_monitor_317;
    df_fifo_intf fifo_intf_318(clock,reset);
    assign fifo_intf_318.rd_en = AESL_inst_myproject.layer2_out_317_U.if_read & AESL_inst_myproject.layer2_out_317_U.if_empty_n;
    assign fifo_intf_318.wr_en = AESL_inst_myproject.layer2_out_317_U.if_write & AESL_inst_myproject.layer2_out_317_U.if_full_n;
    assign fifo_intf_318.fifo_rd_block = 0;
    assign fifo_intf_318.fifo_wr_block = 0;
    assign fifo_intf_318.finish = finish;
    csv_file_dump fifo_csv_dumper_318;
    csv_file_dump cstatus_csv_dumper_318;
    df_fifo_monitor fifo_monitor_318;
    df_fifo_intf fifo_intf_319(clock,reset);
    assign fifo_intf_319.rd_en = AESL_inst_myproject.layer2_out_318_U.if_read & AESL_inst_myproject.layer2_out_318_U.if_empty_n;
    assign fifo_intf_319.wr_en = AESL_inst_myproject.layer2_out_318_U.if_write & AESL_inst_myproject.layer2_out_318_U.if_full_n;
    assign fifo_intf_319.fifo_rd_block = 0;
    assign fifo_intf_319.fifo_wr_block = 0;
    assign fifo_intf_319.finish = finish;
    csv_file_dump fifo_csv_dumper_319;
    csv_file_dump cstatus_csv_dumper_319;
    df_fifo_monitor fifo_monitor_319;
    df_fifo_intf fifo_intf_320(clock,reset);
    assign fifo_intf_320.rd_en = AESL_inst_myproject.layer2_out_319_U.if_read & AESL_inst_myproject.layer2_out_319_U.if_empty_n;
    assign fifo_intf_320.wr_en = AESL_inst_myproject.layer2_out_319_U.if_write & AESL_inst_myproject.layer2_out_319_U.if_full_n;
    assign fifo_intf_320.fifo_rd_block = 0;
    assign fifo_intf_320.fifo_wr_block = 0;
    assign fifo_intf_320.finish = finish;
    csv_file_dump fifo_csv_dumper_320;
    csv_file_dump cstatus_csv_dumper_320;
    df_fifo_monitor fifo_monitor_320;
    df_fifo_intf fifo_intf_321(clock,reset);
    assign fifo_intf_321.rd_en = AESL_inst_myproject.layer2_out_320_U.if_read & AESL_inst_myproject.layer2_out_320_U.if_empty_n;
    assign fifo_intf_321.wr_en = AESL_inst_myproject.layer2_out_320_U.if_write & AESL_inst_myproject.layer2_out_320_U.if_full_n;
    assign fifo_intf_321.fifo_rd_block = 0;
    assign fifo_intf_321.fifo_wr_block = 0;
    assign fifo_intf_321.finish = finish;
    csv_file_dump fifo_csv_dumper_321;
    csv_file_dump cstatus_csv_dumper_321;
    df_fifo_monitor fifo_monitor_321;
    df_fifo_intf fifo_intf_322(clock,reset);
    assign fifo_intf_322.rd_en = AESL_inst_myproject.layer2_out_321_U.if_read & AESL_inst_myproject.layer2_out_321_U.if_empty_n;
    assign fifo_intf_322.wr_en = AESL_inst_myproject.layer2_out_321_U.if_write & AESL_inst_myproject.layer2_out_321_U.if_full_n;
    assign fifo_intf_322.fifo_rd_block = 0;
    assign fifo_intf_322.fifo_wr_block = 0;
    assign fifo_intf_322.finish = finish;
    csv_file_dump fifo_csv_dumper_322;
    csv_file_dump cstatus_csv_dumper_322;
    df_fifo_monitor fifo_monitor_322;
    df_fifo_intf fifo_intf_323(clock,reset);
    assign fifo_intf_323.rd_en = AESL_inst_myproject.layer2_out_322_U.if_read & AESL_inst_myproject.layer2_out_322_U.if_empty_n;
    assign fifo_intf_323.wr_en = AESL_inst_myproject.layer2_out_322_U.if_write & AESL_inst_myproject.layer2_out_322_U.if_full_n;
    assign fifo_intf_323.fifo_rd_block = 0;
    assign fifo_intf_323.fifo_wr_block = 0;
    assign fifo_intf_323.finish = finish;
    csv_file_dump fifo_csv_dumper_323;
    csv_file_dump cstatus_csv_dumper_323;
    df_fifo_monitor fifo_monitor_323;
    df_fifo_intf fifo_intf_324(clock,reset);
    assign fifo_intf_324.rd_en = AESL_inst_myproject.layer2_out_323_U.if_read & AESL_inst_myproject.layer2_out_323_U.if_empty_n;
    assign fifo_intf_324.wr_en = AESL_inst_myproject.layer2_out_323_U.if_write & AESL_inst_myproject.layer2_out_323_U.if_full_n;
    assign fifo_intf_324.fifo_rd_block = 0;
    assign fifo_intf_324.fifo_wr_block = 0;
    assign fifo_intf_324.finish = finish;
    csv_file_dump fifo_csv_dumper_324;
    csv_file_dump cstatus_csv_dumper_324;
    df_fifo_monitor fifo_monitor_324;
    df_fifo_intf fifo_intf_325(clock,reset);
    assign fifo_intf_325.rd_en = AESL_inst_myproject.layer2_out_324_U.if_read & AESL_inst_myproject.layer2_out_324_U.if_empty_n;
    assign fifo_intf_325.wr_en = AESL_inst_myproject.layer2_out_324_U.if_write & AESL_inst_myproject.layer2_out_324_U.if_full_n;
    assign fifo_intf_325.fifo_rd_block = 0;
    assign fifo_intf_325.fifo_wr_block = 0;
    assign fifo_intf_325.finish = finish;
    csv_file_dump fifo_csv_dumper_325;
    csv_file_dump cstatus_csv_dumper_325;
    df_fifo_monitor fifo_monitor_325;
    df_fifo_intf fifo_intf_326(clock,reset);
    assign fifo_intf_326.rd_en = AESL_inst_myproject.layer2_out_325_U.if_read & AESL_inst_myproject.layer2_out_325_U.if_empty_n;
    assign fifo_intf_326.wr_en = AESL_inst_myproject.layer2_out_325_U.if_write & AESL_inst_myproject.layer2_out_325_U.if_full_n;
    assign fifo_intf_326.fifo_rd_block = 0;
    assign fifo_intf_326.fifo_wr_block = 0;
    assign fifo_intf_326.finish = finish;
    csv_file_dump fifo_csv_dumper_326;
    csv_file_dump cstatus_csv_dumper_326;
    df_fifo_monitor fifo_monitor_326;
    df_fifo_intf fifo_intf_327(clock,reset);
    assign fifo_intf_327.rd_en = AESL_inst_myproject.layer2_out_326_U.if_read & AESL_inst_myproject.layer2_out_326_U.if_empty_n;
    assign fifo_intf_327.wr_en = AESL_inst_myproject.layer2_out_326_U.if_write & AESL_inst_myproject.layer2_out_326_U.if_full_n;
    assign fifo_intf_327.fifo_rd_block = 0;
    assign fifo_intf_327.fifo_wr_block = 0;
    assign fifo_intf_327.finish = finish;
    csv_file_dump fifo_csv_dumper_327;
    csv_file_dump cstatus_csv_dumper_327;
    df_fifo_monitor fifo_monitor_327;
    df_fifo_intf fifo_intf_328(clock,reset);
    assign fifo_intf_328.rd_en = AESL_inst_myproject.layer2_out_327_U.if_read & AESL_inst_myproject.layer2_out_327_U.if_empty_n;
    assign fifo_intf_328.wr_en = AESL_inst_myproject.layer2_out_327_U.if_write & AESL_inst_myproject.layer2_out_327_U.if_full_n;
    assign fifo_intf_328.fifo_rd_block = 0;
    assign fifo_intf_328.fifo_wr_block = 0;
    assign fifo_intf_328.finish = finish;
    csv_file_dump fifo_csv_dumper_328;
    csv_file_dump cstatus_csv_dumper_328;
    df_fifo_monitor fifo_monitor_328;
    df_fifo_intf fifo_intf_329(clock,reset);
    assign fifo_intf_329.rd_en = AESL_inst_myproject.layer2_out_328_U.if_read & AESL_inst_myproject.layer2_out_328_U.if_empty_n;
    assign fifo_intf_329.wr_en = AESL_inst_myproject.layer2_out_328_U.if_write & AESL_inst_myproject.layer2_out_328_U.if_full_n;
    assign fifo_intf_329.fifo_rd_block = 0;
    assign fifo_intf_329.fifo_wr_block = 0;
    assign fifo_intf_329.finish = finish;
    csv_file_dump fifo_csv_dumper_329;
    csv_file_dump cstatus_csv_dumper_329;
    df_fifo_monitor fifo_monitor_329;
    df_fifo_intf fifo_intf_330(clock,reset);
    assign fifo_intf_330.rd_en = AESL_inst_myproject.layer2_out_329_U.if_read & AESL_inst_myproject.layer2_out_329_U.if_empty_n;
    assign fifo_intf_330.wr_en = AESL_inst_myproject.layer2_out_329_U.if_write & AESL_inst_myproject.layer2_out_329_U.if_full_n;
    assign fifo_intf_330.fifo_rd_block = 0;
    assign fifo_intf_330.fifo_wr_block = 0;
    assign fifo_intf_330.finish = finish;
    csv_file_dump fifo_csv_dumper_330;
    csv_file_dump cstatus_csv_dumper_330;
    df_fifo_monitor fifo_monitor_330;
    df_fifo_intf fifo_intf_331(clock,reset);
    assign fifo_intf_331.rd_en = AESL_inst_myproject.layer2_out_330_U.if_read & AESL_inst_myproject.layer2_out_330_U.if_empty_n;
    assign fifo_intf_331.wr_en = AESL_inst_myproject.layer2_out_330_U.if_write & AESL_inst_myproject.layer2_out_330_U.if_full_n;
    assign fifo_intf_331.fifo_rd_block = 0;
    assign fifo_intf_331.fifo_wr_block = 0;
    assign fifo_intf_331.finish = finish;
    csv_file_dump fifo_csv_dumper_331;
    csv_file_dump cstatus_csv_dumper_331;
    df_fifo_monitor fifo_monitor_331;
    df_fifo_intf fifo_intf_332(clock,reset);
    assign fifo_intf_332.rd_en = AESL_inst_myproject.layer2_out_331_U.if_read & AESL_inst_myproject.layer2_out_331_U.if_empty_n;
    assign fifo_intf_332.wr_en = AESL_inst_myproject.layer2_out_331_U.if_write & AESL_inst_myproject.layer2_out_331_U.if_full_n;
    assign fifo_intf_332.fifo_rd_block = 0;
    assign fifo_intf_332.fifo_wr_block = 0;
    assign fifo_intf_332.finish = finish;
    csv_file_dump fifo_csv_dumper_332;
    csv_file_dump cstatus_csv_dumper_332;
    df_fifo_monitor fifo_monitor_332;
    df_fifo_intf fifo_intf_333(clock,reset);
    assign fifo_intf_333.rd_en = AESL_inst_myproject.layer2_out_332_U.if_read & AESL_inst_myproject.layer2_out_332_U.if_empty_n;
    assign fifo_intf_333.wr_en = AESL_inst_myproject.layer2_out_332_U.if_write & AESL_inst_myproject.layer2_out_332_U.if_full_n;
    assign fifo_intf_333.fifo_rd_block = 0;
    assign fifo_intf_333.fifo_wr_block = 0;
    assign fifo_intf_333.finish = finish;
    csv_file_dump fifo_csv_dumper_333;
    csv_file_dump cstatus_csv_dumper_333;
    df_fifo_monitor fifo_monitor_333;
    df_fifo_intf fifo_intf_334(clock,reset);
    assign fifo_intf_334.rd_en = AESL_inst_myproject.layer2_out_333_U.if_read & AESL_inst_myproject.layer2_out_333_U.if_empty_n;
    assign fifo_intf_334.wr_en = AESL_inst_myproject.layer2_out_333_U.if_write & AESL_inst_myproject.layer2_out_333_U.if_full_n;
    assign fifo_intf_334.fifo_rd_block = 0;
    assign fifo_intf_334.fifo_wr_block = 0;
    assign fifo_intf_334.finish = finish;
    csv_file_dump fifo_csv_dumper_334;
    csv_file_dump cstatus_csv_dumper_334;
    df_fifo_monitor fifo_monitor_334;
    df_fifo_intf fifo_intf_335(clock,reset);
    assign fifo_intf_335.rd_en = AESL_inst_myproject.layer2_out_334_U.if_read & AESL_inst_myproject.layer2_out_334_U.if_empty_n;
    assign fifo_intf_335.wr_en = AESL_inst_myproject.layer2_out_334_U.if_write & AESL_inst_myproject.layer2_out_334_U.if_full_n;
    assign fifo_intf_335.fifo_rd_block = 0;
    assign fifo_intf_335.fifo_wr_block = 0;
    assign fifo_intf_335.finish = finish;
    csv_file_dump fifo_csv_dumper_335;
    csv_file_dump cstatus_csv_dumper_335;
    df_fifo_monitor fifo_monitor_335;
    df_fifo_intf fifo_intf_336(clock,reset);
    assign fifo_intf_336.rd_en = AESL_inst_myproject.layer2_out_335_U.if_read & AESL_inst_myproject.layer2_out_335_U.if_empty_n;
    assign fifo_intf_336.wr_en = AESL_inst_myproject.layer2_out_335_U.if_write & AESL_inst_myproject.layer2_out_335_U.if_full_n;
    assign fifo_intf_336.fifo_rd_block = 0;
    assign fifo_intf_336.fifo_wr_block = 0;
    assign fifo_intf_336.finish = finish;
    csv_file_dump fifo_csv_dumper_336;
    csv_file_dump cstatus_csv_dumper_336;
    df_fifo_monitor fifo_monitor_336;
    df_fifo_intf fifo_intf_337(clock,reset);
    assign fifo_intf_337.rd_en = AESL_inst_myproject.layer2_out_336_U.if_read & AESL_inst_myproject.layer2_out_336_U.if_empty_n;
    assign fifo_intf_337.wr_en = AESL_inst_myproject.layer2_out_336_U.if_write & AESL_inst_myproject.layer2_out_336_U.if_full_n;
    assign fifo_intf_337.fifo_rd_block = 0;
    assign fifo_intf_337.fifo_wr_block = 0;
    assign fifo_intf_337.finish = finish;
    csv_file_dump fifo_csv_dumper_337;
    csv_file_dump cstatus_csv_dumper_337;
    df_fifo_monitor fifo_monitor_337;
    df_fifo_intf fifo_intf_338(clock,reset);
    assign fifo_intf_338.rd_en = AESL_inst_myproject.layer2_out_337_U.if_read & AESL_inst_myproject.layer2_out_337_U.if_empty_n;
    assign fifo_intf_338.wr_en = AESL_inst_myproject.layer2_out_337_U.if_write & AESL_inst_myproject.layer2_out_337_U.if_full_n;
    assign fifo_intf_338.fifo_rd_block = 0;
    assign fifo_intf_338.fifo_wr_block = 0;
    assign fifo_intf_338.finish = finish;
    csv_file_dump fifo_csv_dumper_338;
    csv_file_dump cstatus_csv_dumper_338;
    df_fifo_monitor fifo_monitor_338;
    df_fifo_intf fifo_intf_339(clock,reset);
    assign fifo_intf_339.rd_en = AESL_inst_myproject.layer2_out_338_U.if_read & AESL_inst_myproject.layer2_out_338_U.if_empty_n;
    assign fifo_intf_339.wr_en = AESL_inst_myproject.layer2_out_338_U.if_write & AESL_inst_myproject.layer2_out_338_U.if_full_n;
    assign fifo_intf_339.fifo_rd_block = 0;
    assign fifo_intf_339.fifo_wr_block = 0;
    assign fifo_intf_339.finish = finish;
    csv_file_dump fifo_csv_dumper_339;
    csv_file_dump cstatus_csv_dumper_339;
    df_fifo_monitor fifo_monitor_339;
    df_fifo_intf fifo_intf_340(clock,reset);
    assign fifo_intf_340.rd_en = AESL_inst_myproject.layer2_out_339_U.if_read & AESL_inst_myproject.layer2_out_339_U.if_empty_n;
    assign fifo_intf_340.wr_en = AESL_inst_myproject.layer2_out_339_U.if_write & AESL_inst_myproject.layer2_out_339_U.if_full_n;
    assign fifo_intf_340.fifo_rd_block = 0;
    assign fifo_intf_340.fifo_wr_block = 0;
    assign fifo_intf_340.finish = finish;
    csv_file_dump fifo_csv_dumper_340;
    csv_file_dump cstatus_csv_dumper_340;
    df_fifo_monitor fifo_monitor_340;
    df_fifo_intf fifo_intf_341(clock,reset);
    assign fifo_intf_341.rd_en = AESL_inst_myproject.layer2_out_340_U.if_read & AESL_inst_myproject.layer2_out_340_U.if_empty_n;
    assign fifo_intf_341.wr_en = AESL_inst_myproject.layer2_out_340_U.if_write & AESL_inst_myproject.layer2_out_340_U.if_full_n;
    assign fifo_intf_341.fifo_rd_block = 0;
    assign fifo_intf_341.fifo_wr_block = 0;
    assign fifo_intf_341.finish = finish;
    csv_file_dump fifo_csv_dumper_341;
    csv_file_dump cstatus_csv_dumper_341;
    df_fifo_monitor fifo_monitor_341;
    df_fifo_intf fifo_intf_342(clock,reset);
    assign fifo_intf_342.rd_en = AESL_inst_myproject.layer2_out_341_U.if_read & AESL_inst_myproject.layer2_out_341_U.if_empty_n;
    assign fifo_intf_342.wr_en = AESL_inst_myproject.layer2_out_341_U.if_write & AESL_inst_myproject.layer2_out_341_U.if_full_n;
    assign fifo_intf_342.fifo_rd_block = 0;
    assign fifo_intf_342.fifo_wr_block = 0;
    assign fifo_intf_342.finish = finish;
    csv_file_dump fifo_csv_dumper_342;
    csv_file_dump cstatus_csv_dumper_342;
    df_fifo_monitor fifo_monitor_342;
    df_fifo_intf fifo_intf_343(clock,reset);
    assign fifo_intf_343.rd_en = AESL_inst_myproject.layer2_out_342_U.if_read & AESL_inst_myproject.layer2_out_342_U.if_empty_n;
    assign fifo_intf_343.wr_en = AESL_inst_myproject.layer2_out_342_U.if_write & AESL_inst_myproject.layer2_out_342_U.if_full_n;
    assign fifo_intf_343.fifo_rd_block = 0;
    assign fifo_intf_343.fifo_wr_block = 0;
    assign fifo_intf_343.finish = finish;
    csv_file_dump fifo_csv_dumper_343;
    csv_file_dump cstatus_csv_dumper_343;
    df_fifo_monitor fifo_monitor_343;
    df_fifo_intf fifo_intf_344(clock,reset);
    assign fifo_intf_344.rd_en = AESL_inst_myproject.layer2_out_343_U.if_read & AESL_inst_myproject.layer2_out_343_U.if_empty_n;
    assign fifo_intf_344.wr_en = AESL_inst_myproject.layer2_out_343_U.if_write & AESL_inst_myproject.layer2_out_343_U.if_full_n;
    assign fifo_intf_344.fifo_rd_block = 0;
    assign fifo_intf_344.fifo_wr_block = 0;
    assign fifo_intf_344.finish = finish;
    csv_file_dump fifo_csv_dumper_344;
    csv_file_dump cstatus_csv_dumper_344;
    df_fifo_monitor fifo_monitor_344;
    df_fifo_intf fifo_intf_345(clock,reset);
    assign fifo_intf_345.rd_en = AESL_inst_myproject.layer2_out_344_U.if_read & AESL_inst_myproject.layer2_out_344_U.if_empty_n;
    assign fifo_intf_345.wr_en = AESL_inst_myproject.layer2_out_344_U.if_write & AESL_inst_myproject.layer2_out_344_U.if_full_n;
    assign fifo_intf_345.fifo_rd_block = 0;
    assign fifo_intf_345.fifo_wr_block = 0;
    assign fifo_intf_345.finish = finish;
    csv_file_dump fifo_csv_dumper_345;
    csv_file_dump cstatus_csv_dumper_345;
    df_fifo_monitor fifo_monitor_345;
    df_fifo_intf fifo_intf_346(clock,reset);
    assign fifo_intf_346.rd_en = AESL_inst_myproject.layer2_out_345_U.if_read & AESL_inst_myproject.layer2_out_345_U.if_empty_n;
    assign fifo_intf_346.wr_en = AESL_inst_myproject.layer2_out_345_U.if_write & AESL_inst_myproject.layer2_out_345_U.if_full_n;
    assign fifo_intf_346.fifo_rd_block = 0;
    assign fifo_intf_346.fifo_wr_block = 0;
    assign fifo_intf_346.finish = finish;
    csv_file_dump fifo_csv_dumper_346;
    csv_file_dump cstatus_csv_dumper_346;
    df_fifo_monitor fifo_monitor_346;
    df_fifo_intf fifo_intf_347(clock,reset);
    assign fifo_intf_347.rd_en = AESL_inst_myproject.layer2_out_346_U.if_read & AESL_inst_myproject.layer2_out_346_U.if_empty_n;
    assign fifo_intf_347.wr_en = AESL_inst_myproject.layer2_out_346_U.if_write & AESL_inst_myproject.layer2_out_346_U.if_full_n;
    assign fifo_intf_347.fifo_rd_block = 0;
    assign fifo_intf_347.fifo_wr_block = 0;
    assign fifo_intf_347.finish = finish;
    csv_file_dump fifo_csv_dumper_347;
    csv_file_dump cstatus_csv_dumper_347;
    df_fifo_monitor fifo_monitor_347;
    df_fifo_intf fifo_intf_348(clock,reset);
    assign fifo_intf_348.rd_en = AESL_inst_myproject.layer2_out_347_U.if_read & AESL_inst_myproject.layer2_out_347_U.if_empty_n;
    assign fifo_intf_348.wr_en = AESL_inst_myproject.layer2_out_347_U.if_write & AESL_inst_myproject.layer2_out_347_U.if_full_n;
    assign fifo_intf_348.fifo_rd_block = 0;
    assign fifo_intf_348.fifo_wr_block = 0;
    assign fifo_intf_348.finish = finish;
    csv_file_dump fifo_csv_dumper_348;
    csv_file_dump cstatus_csv_dumper_348;
    df_fifo_monitor fifo_monitor_348;
    df_fifo_intf fifo_intf_349(clock,reset);
    assign fifo_intf_349.rd_en = AESL_inst_myproject.layer2_out_348_U.if_read & AESL_inst_myproject.layer2_out_348_U.if_empty_n;
    assign fifo_intf_349.wr_en = AESL_inst_myproject.layer2_out_348_U.if_write & AESL_inst_myproject.layer2_out_348_U.if_full_n;
    assign fifo_intf_349.fifo_rd_block = 0;
    assign fifo_intf_349.fifo_wr_block = 0;
    assign fifo_intf_349.finish = finish;
    csv_file_dump fifo_csv_dumper_349;
    csv_file_dump cstatus_csv_dumper_349;
    df_fifo_monitor fifo_monitor_349;
    df_fifo_intf fifo_intf_350(clock,reset);
    assign fifo_intf_350.rd_en = AESL_inst_myproject.layer2_out_349_U.if_read & AESL_inst_myproject.layer2_out_349_U.if_empty_n;
    assign fifo_intf_350.wr_en = AESL_inst_myproject.layer2_out_349_U.if_write & AESL_inst_myproject.layer2_out_349_U.if_full_n;
    assign fifo_intf_350.fifo_rd_block = 0;
    assign fifo_intf_350.fifo_wr_block = 0;
    assign fifo_intf_350.finish = finish;
    csv_file_dump fifo_csv_dumper_350;
    csv_file_dump cstatus_csv_dumper_350;
    df_fifo_monitor fifo_monitor_350;
    df_fifo_intf fifo_intf_351(clock,reset);
    assign fifo_intf_351.rd_en = AESL_inst_myproject.layer2_out_350_U.if_read & AESL_inst_myproject.layer2_out_350_U.if_empty_n;
    assign fifo_intf_351.wr_en = AESL_inst_myproject.layer2_out_350_U.if_write & AESL_inst_myproject.layer2_out_350_U.if_full_n;
    assign fifo_intf_351.fifo_rd_block = 0;
    assign fifo_intf_351.fifo_wr_block = 0;
    assign fifo_intf_351.finish = finish;
    csv_file_dump fifo_csv_dumper_351;
    csv_file_dump cstatus_csv_dumper_351;
    df_fifo_monitor fifo_monitor_351;
    df_fifo_intf fifo_intf_352(clock,reset);
    assign fifo_intf_352.rd_en = AESL_inst_myproject.layer2_out_351_U.if_read & AESL_inst_myproject.layer2_out_351_U.if_empty_n;
    assign fifo_intf_352.wr_en = AESL_inst_myproject.layer2_out_351_U.if_write & AESL_inst_myproject.layer2_out_351_U.if_full_n;
    assign fifo_intf_352.fifo_rd_block = 0;
    assign fifo_intf_352.fifo_wr_block = 0;
    assign fifo_intf_352.finish = finish;
    csv_file_dump fifo_csv_dumper_352;
    csv_file_dump cstatus_csv_dumper_352;
    df_fifo_monitor fifo_monitor_352;
    df_fifo_intf fifo_intf_353(clock,reset);
    assign fifo_intf_353.rd_en = AESL_inst_myproject.layer2_out_352_U.if_read & AESL_inst_myproject.layer2_out_352_U.if_empty_n;
    assign fifo_intf_353.wr_en = AESL_inst_myproject.layer2_out_352_U.if_write & AESL_inst_myproject.layer2_out_352_U.if_full_n;
    assign fifo_intf_353.fifo_rd_block = 0;
    assign fifo_intf_353.fifo_wr_block = 0;
    assign fifo_intf_353.finish = finish;
    csv_file_dump fifo_csv_dumper_353;
    csv_file_dump cstatus_csv_dumper_353;
    df_fifo_monitor fifo_monitor_353;
    df_fifo_intf fifo_intf_354(clock,reset);
    assign fifo_intf_354.rd_en = AESL_inst_myproject.layer2_out_353_U.if_read & AESL_inst_myproject.layer2_out_353_U.if_empty_n;
    assign fifo_intf_354.wr_en = AESL_inst_myproject.layer2_out_353_U.if_write & AESL_inst_myproject.layer2_out_353_U.if_full_n;
    assign fifo_intf_354.fifo_rd_block = 0;
    assign fifo_intf_354.fifo_wr_block = 0;
    assign fifo_intf_354.finish = finish;
    csv_file_dump fifo_csv_dumper_354;
    csv_file_dump cstatus_csv_dumper_354;
    df_fifo_monitor fifo_monitor_354;
    df_fifo_intf fifo_intf_355(clock,reset);
    assign fifo_intf_355.rd_en = AESL_inst_myproject.layer2_out_354_U.if_read & AESL_inst_myproject.layer2_out_354_U.if_empty_n;
    assign fifo_intf_355.wr_en = AESL_inst_myproject.layer2_out_354_U.if_write & AESL_inst_myproject.layer2_out_354_U.if_full_n;
    assign fifo_intf_355.fifo_rd_block = 0;
    assign fifo_intf_355.fifo_wr_block = 0;
    assign fifo_intf_355.finish = finish;
    csv_file_dump fifo_csv_dumper_355;
    csv_file_dump cstatus_csv_dumper_355;
    df_fifo_monitor fifo_monitor_355;
    df_fifo_intf fifo_intf_356(clock,reset);
    assign fifo_intf_356.rd_en = AESL_inst_myproject.layer2_out_355_U.if_read & AESL_inst_myproject.layer2_out_355_U.if_empty_n;
    assign fifo_intf_356.wr_en = AESL_inst_myproject.layer2_out_355_U.if_write & AESL_inst_myproject.layer2_out_355_U.if_full_n;
    assign fifo_intf_356.fifo_rd_block = 0;
    assign fifo_intf_356.fifo_wr_block = 0;
    assign fifo_intf_356.finish = finish;
    csv_file_dump fifo_csv_dumper_356;
    csv_file_dump cstatus_csv_dumper_356;
    df_fifo_monitor fifo_monitor_356;
    df_fifo_intf fifo_intf_357(clock,reset);
    assign fifo_intf_357.rd_en = AESL_inst_myproject.layer2_out_356_U.if_read & AESL_inst_myproject.layer2_out_356_U.if_empty_n;
    assign fifo_intf_357.wr_en = AESL_inst_myproject.layer2_out_356_U.if_write & AESL_inst_myproject.layer2_out_356_U.if_full_n;
    assign fifo_intf_357.fifo_rd_block = 0;
    assign fifo_intf_357.fifo_wr_block = 0;
    assign fifo_intf_357.finish = finish;
    csv_file_dump fifo_csv_dumper_357;
    csv_file_dump cstatus_csv_dumper_357;
    df_fifo_monitor fifo_monitor_357;
    df_fifo_intf fifo_intf_358(clock,reset);
    assign fifo_intf_358.rd_en = AESL_inst_myproject.layer2_out_357_U.if_read & AESL_inst_myproject.layer2_out_357_U.if_empty_n;
    assign fifo_intf_358.wr_en = AESL_inst_myproject.layer2_out_357_U.if_write & AESL_inst_myproject.layer2_out_357_U.if_full_n;
    assign fifo_intf_358.fifo_rd_block = 0;
    assign fifo_intf_358.fifo_wr_block = 0;
    assign fifo_intf_358.finish = finish;
    csv_file_dump fifo_csv_dumper_358;
    csv_file_dump cstatus_csv_dumper_358;
    df_fifo_monitor fifo_monitor_358;
    df_fifo_intf fifo_intf_359(clock,reset);
    assign fifo_intf_359.rd_en = AESL_inst_myproject.layer2_out_358_U.if_read & AESL_inst_myproject.layer2_out_358_U.if_empty_n;
    assign fifo_intf_359.wr_en = AESL_inst_myproject.layer2_out_358_U.if_write & AESL_inst_myproject.layer2_out_358_U.if_full_n;
    assign fifo_intf_359.fifo_rd_block = 0;
    assign fifo_intf_359.fifo_wr_block = 0;
    assign fifo_intf_359.finish = finish;
    csv_file_dump fifo_csv_dumper_359;
    csv_file_dump cstatus_csv_dumper_359;
    df_fifo_monitor fifo_monitor_359;
    df_fifo_intf fifo_intf_360(clock,reset);
    assign fifo_intf_360.rd_en = AESL_inst_myproject.layer2_out_359_U.if_read & AESL_inst_myproject.layer2_out_359_U.if_empty_n;
    assign fifo_intf_360.wr_en = AESL_inst_myproject.layer2_out_359_U.if_write & AESL_inst_myproject.layer2_out_359_U.if_full_n;
    assign fifo_intf_360.fifo_rd_block = 0;
    assign fifo_intf_360.fifo_wr_block = 0;
    assign fifo_intf_360.finish = finish;
    csv_file_dump fifo_csv_dumper_360;
    csv_file_dump cstatus_csv_dumper_360;
    df_fifo_monitor fifo_monitor_360;
    df_fifo_intf fifo_intf_361(clock,reset);
    assign fifo_intf_361.rd_en = AESL_inst_myproject.layer2_out_360_U.if_read & AESL_inst_myproject.layer2_out_360_U.if_empty_n;
    assign fifo_intf_361.wr_en = AESL_inst_myproject.layer2_out_360_U.if_write & AESL_inst_myproject.layer2_out_360_U.if_full_n;
    assign fifo_intf_361.fifo_rd_block = 0;
    assign fifo_intf_361.fifo_wr_block = 0;
    assign fifo_intf_361.finish = finish;
    csv_file_dump fifo_csv_dumper_361;
    csv_file_dump cstatus_csv_dumper_361;
    df_fifo_monitor fifo_monitor_361;
    df_fifo_intf fifo_intf_362(clock,reset);
    assign fifo_intf_362.rd_en = AESL_inst_myproject.layer2_out_361_U.if_read & AESL_inst_myproject.layer2_out_361_U.if_empty_n;
    assign fifo_intf_362.wr_en = AESL_inst_myproject.layer2_out_361_U.if_write & AESL_inst_myproject.layer2_out_361_U.if_full_n;
    assign fifo_intf_362.fifo_rd_block = 0;
    assign fifo_intf_362.fifo_wr_block = 0;
    assign fifo_intf_362.finish = finish;
    csv_file_dump fifo_csv_dumper_362;
    csv_file_dump cstatus_csv_dumper_362;
    df_fifo_monitor fifo_monitor_362;
    df_fifo_intf fifo_intf_363(clock,reset);
    assign fifo_intf_363.rd_en = AESL_inst_myproject.layer2_out_362_U.if_read & AESL_inst_myproject.layer2_out_362_U.if_empty_n;
    assign fifo_intf_363.wr_en = AESL_inst_myproject.layer2_out_362_U.if_write & AESL_inst_myproject.layer2_out_362_U.if_full_n;
    assign fifo_intf_363.fifo_rd_block = 0;
    assign fifo_intf_363.fifo_wr_block = 0;
    assign fifo_intf_363.finish = finish;
    csv_file_dump fifo_csv_dumper_363;
    csv_file_dump cstatus_csv_dumper_363;
    df_fifo_monitor fifo_monitor_363;
    df_fifo_intf fifo_intf_364(clock,reset);
    assign fifo_intf_364.rd_en = AESL_inst_myproject.layer2_out_363_U.if_read & AESL_inst_myproject.layer2_out_363_U.if_empty_n;
    assign fifo_intf_364.wr_en = AESL_inst_myproject.layer2_out_363_U.if_write & AESL_inst_myproject.layer2_out_363_U.if_full_n;
    assign fifo_intf_364.fifo_rd_block = 0;
    assign fifo_intf_364.fifo_wr_block = 0;
    assign fifo_intf_364.finish = finish;
    csv_file_dump fifo_csv_dumper_364;
    csv_file_dump cstatus_csv_dumper_364;
    df_fifo_monitor fifo_monitor_364;
    df_fifo_intf fifo_intf_365(clock,reset);
    assign fifo_intf_365.rd_en = AESL_inst_myproject.layer2_out_364_U.if_read & AESL_inst_myproject.layer2_out_364_U.if_empty_n;
    assign fifo_intf_365.wr_en = AESL_inst_myproject.layer2_out_364_U.if_write & AESL_inst_myproject.layer2_out_364_U.if_full_n;
    assign fifo_intf_365.fifo_rd_block = 0;
    assign fifo_intf_365.fifo_wr_block = 0;
    assign fifo_intf_365.finish = finish;
    csv_file_dump fifo_csv_dumper_365;
    csv_file_dump cstatus_csv_dumper_365;
    df_fifo_monitor fifo_monitor_365;
    df_fifo_intf fifo_intf_366(clock,reset);
    assign fifo_intf_366.rd_en = AESL_inst_myproject.layer2_out_365_U.if_read & AESL_inst_myproject.layer2_out_365_U.if_empty_n;
    assign fifo_intf_366.wr_en = AESL_inst_myproject.layer2_out_365_U.if_write & AESL_inst_myproject.layer2_out_365_U.if_full_n;
    assign fifo_intf_366.fifo_rd_block = 0;
    assign fifo_intf_366.fifo_wr_block = 0;
    assign fifo_intf_366.finish = finish;
    csv_file_dump fifo_csv_dumper_366;
    csv_file_dump cstatus_csv_dumper_366;
    df_fifo_monitor fifo_monitor_366;
    df_fifo_intf fifo_intf_367(clock,reset);
    assign fifo_intf_367.rd_en = AESL_inst_myproject.layer2_out_366_U.if_read & AESL_inst_myproject.layer2_out_366_U.if_empty_n;
    assign fifo_intf_367.wr_en = AESL_inst_myproject.layer2_out_366_U.if_write & AESL_inst_myproject.layer2_out_366_U.if_full_n;
    assign fifo_intf_367.fifo_rd_block = 0;
    assign fifo_intf_367.fifo_wr_block = 0;
    assign fifo_intf_367.finish = finish;
    csv_file_dump fifo_csv_dumper_367;
    csv_file_dump cstatus_csv_dumper_367;
    df_fifo_monitor fifo_monitor_367;
    df_fifo_intf fifo_intf_368(clock,reset);
    assign fifo_intf_368.rd_en = AESL_inst_myproject.layer2_out_367_U.if_read & AESL_inst_myproject.layer2_out_367_U.if_empty_n;
    assign fifo_intf_368.wr_en = AESL_inst_myproject.layer2_out_367_U.if_write & AESL_inst_myproject.layer2_out_367_U.if_full_n;
    assign fifo_intf_368.fifo_rd_block = 0;
    assign fifo_intf_368.fifo_wr_block = 0;
    assign fifo_intf_368.finish = finish;
    csv_file_dump fifo_csv_dumper_368;
    csv_file_dump cstatus_csv_dumper_368;
    df_fifo_monitor fifo_monitor_368;
    df_fifo_intf fifo_intf_369(clock,reset);
    assign fifo_intf_369.rd_en = AESL_inst_myproject.layer2_out_368_U.if_read & AESL_inst_myproject.layer2_out_368_U.if_empty_n;
    assign fifo_intf_369.wr_en = AESL_inst_myproject.layer2_out_368_U.if_write & AESL_inst_myproject.layer2_out_368_U.if_full_n;
    assign fifo_intf_369.fifo_rd_block = 0;
    assign fifo_intf_369.fifo_wr_block = 0;
    assign fifo_intf_369.finish = finish;
    csv_file_dump fifo_csv_dumper_369;
    csv_file_dump cstatus_csv_dumper_369;
    df_fifo_monitor fifo_monitor_369;
    df_fifo_intf fifo_intf_370(clock,reset);
    assign fifo_intf_370.rd_en = AESL_inst_myproject.layer2_out_369_U.if_read & AESL_inst_myproject.layer2_out_369_U.if_empty_n;
    assign fifo_intf_370.wr_en = AESL_inst_myproject.layer2_out_369_U.if_write & AESL_inst_myproject.layer2_out_369_U.if_full_n;
    assign fifo_intf_370.fifo_rd_block = 0;
    assign fifo_intf_370.fifo_wr_block = 0;
    assign fifo_intf_370.finish = finish;
    csv_file_dump fifo_csv_dumper_370;
    csv_file_dump cstatus_csv_dumper_370;
    df_fifo_monitor fifo_monitor_370;
    df_fifo_intf fifo_intf_371(clock,reset);
    assign fifo_intf_371.rd_en = AESL_inst_myproject.layer2_out_370_U.if_read & AESL_inst_myproject.layer2_out_370_U.if_empty_n;
    assign fifo_intf_371.wr_en = AESL_inst_myproject.layer2_out_370_U.if_write & AESL_inst_myproject.layer2_out_370_U.if_full_n;
    assign fifo_intf_371.fifo_rd_block = 0;
    assign fifo_intf_371.fifo_wr_block = 0;
    assign fifo_intf_371.finish = finish;
    csv_file_dump fifo_csv_dumper_371;
    csv_file_dump cstatus_csv_dumper_371;
    df_fifo_monitor fifo_monitor_371;
    df_fifo_intf fifo_intf_372(clock,reset);
    assign fifo_intf_372.rd_en = AESL_inst_myproject.layer2_out_371_U.if_read & AESL_inst_myproject.layer2_out_371_U.if_empty_n;
    assign fifo_intf_372.wr_en = AESL_inst_myproject.layer2_out_371_U.if_write & AESL_inst_myproject.layer2_out_371_U.if_full_n;
    assign fifo_intf_372.fifo_rd_block = 0;
    assign fifo_intf_372.fifo_wr_block = 0;
    assign fifo_intf_372.finish = finish;
    csv_file_dump fifo_csv_dumper_372;
    csv_file_dump cstatus_csv_dumper_372;
    df_fifo_monitor fifo_monitor_372;
    df_fifo_intf fifo_intf_373(clock,reset);
    assign fifo_intf_373.rd_en = AESL_inst_myproject.layer2_out_372_U.if_read & AESL_inst_myproject.layer2_out_372_U.if_empty_n;
    assign fifo_intf_373.wr_en = AESL_inst_myproject.layer2_out_372_U.if_write & AESL_inst_myproject.layer2_out_372_U.if_full_n;
    assign fifo_intf_373.fifo_rd_block = 0;
    assign fifo_intf_373.fifo_wr_block = 0;
    assign fifo_intf_373.finish = finish;
    csv_file_dump fifo_csv_dumper_373;
    csv_file_dump cstatus_csv_dumper_373;
    df_fifo_monitor fifo_monitor_373;
    df_fifo_intf fifo_intf_374(clock,reset);
    assign fifo_intf_374.rd_en = AESL_inst_myproject.layer2_out_373_U.if_read & AESL_inst_myproject.layer2_out_373_U.if_empty_n;
    assign fifo_intf_374.wr_en = AESL_inst_myproject.layer2_out_373_U.if_write & AESL_inst_myproject.layer2_out_373_U.if_full_n;
    assign fifo_intf_374.fifo_rd_block = 0;
    assign fifo_intf_374.fifo_wr_block = 0;
    assign fifo_intf_374.finish = finish;
    csv_file_dump fifo_csv_dumper_374;
    csv_file_dump cstatus_csv_dumper_374;
    df_fifo_monitor fifo_monitor_374;
    df_fifo_intf fifo_intf_375(clock,reset);
    assign fifo_intf_375.rd_en = AESL_inst_myproject.layer2_out_374_U.if_read & AESL_inst_myproject.layer2_out_374_U.if_empty_n;
    assign fifo_intf_375.wr_en = AESL_inst_myproject.layer2_out_374_U.if_write & AESL_inst_myproject.layer2_out_374_U.if_full_n;
    assign fifo_intf_375.fifo_rd_block = 0;
    assign fifo_intf_375.fifo_wr_block = 0;
    assign fifo_intf_375.finish = finish;
    csv_file_dump fifo_csv_dumper_375;
    csv_file_dump cstatus_csv_dumper_375;
    df_fifo_monitor fifo_monitor_375;
    df_fifo_intf fifo_intf_376(clock,reset);
    assign fifo_intf_376.rd_en = AESL_inst_myproject.layer2_out_375_U.if_read & AESL_inst_myproject.layer2_out_375_U.if_empty_n;
    assign fifo_intf_376.wr_en = AESL_inst_myproject.layer2_out_375_U.if_write & AESL_inst_myproject.layer2_out_375_U.if_full_n;
    assign fifo_intf_376.fifo_rd_block = 0;
    assign fifo_intf_376.fifo_wr_block = 0;
    assign fifo_intf_376.finish = finish;
    csv_file_dump fifo_csv_dumper_376;
    csv_file_dump cstatus_csv_dumper_376;
    df_fifo_monitor fifo_monitor_376;
    df_fifo_intf fifo_intf_377(clock,reset);
    assign fifo_intf_377.rd_en = AESL_inst_myproject.layer2_out_376_U.if_read & AESL_inst_myproject.layer2_out_376_U.if_empty_n;
    assign fifo_intf_377.wr_en = AESL_inst_myproject.layer2_out_376_U.if_write & AESL_inst_myproject.layer2_out_376_U.if_full_n;
    assign fifo_intf_377.fifo_rd_block = 0;
    assign fifo_intf_377.fifo_wr_block = 0;
    assign fifo_intf_377.finish = finish;
    csv_file_dump fifo_csv_dumper_377;
    csv_file_dump cstatus_csv_dumper_377;
    df_fifo_monitor fifo_monitor_377;
    df_fifo_intf fifo_intf_378(clock,reset);
    assign fifo_intf_378.rd_en = AESL_inst_myproject.layer2_out_377_U.if_read & AESL_inst_myproject.layer2_out_377_U.if_empty_n;
    assign fifo_intf_378.wr_en = AESL_inst_myproject.layer2_out_377_U.if_write & AESL_inst_myproject.layer2_out_377_U.if_full_n;
    assign fifo_intf_378.fifo_rd_block = 0;
    assign fifo_intf_378.fifo_wr_block = 0;
    assign fifo_intf_378.finish = finish;
    csv_file_dump fifo_csv_dumper_378;
    csv_file_dump cstatus_csv_dumper_378;
    df_fifo_monitor fifo_monitor_378;
    df_fifo_intf fifo_intf_379(clock,reset);
    assign fifo_intf_379.rd_en = AESL_inst_myproject.layer2_out_378_U.if_read & AESL_inst_myproject.layer2_out_378_U.if_empty_n;
    assign fifo_intf_379.wr_en = AESL_inst_myproject.layer2_out_378_U.if_write & AESL_inst_myproject.layer2_out_378_U.if_full_n;
    assign fifo_intf_379.fifo_rd_block = 0;
    assign fifo_intf_379.fifo_wr_block = 0;
    assign fifo_intf_379.finish = finish;
    csv_file_dump fifo_csv_dumper_379;
    csv_file_dump cstatus_csv_dumper_379;
    df_fifo_monitor fifo_monitor_379;
    df_fifo_intf fifo_intf_380(clock,reset);
    assign fifo_intf_380.rd_en = AESL_inst_myproject.layer2_out_379_U.if_read & AESL_inst_myproject.layer2_out_379_U.if_empty_n;
    assign fifo_intf_380.wr_en = AESL_inst_myproject.layer2_out_379_U.if_write & AESL_inst_myproject.layer2_out_379_U.if_full_n;
    assign fifo_intf_380.fifo_rd_block = 0;
    assign fifo_intf_380.fifo_wr_block = 0;
    assign fifo_intf_380.finish = finish;
    csv_file_dump fifo_csv_dumper_380;
    csv_file_dump cstatus_csv_dumper_380;
    df_fifo_monitor fifo_monitor_380;
    df_fifo_intf fifo_intf_381(clock,reset);
    assign fifo_intf_381.rd_en = AESL_inst_myproject.layer2_out_380_U.if_read & AESL_inst_myproject.layer2_out_380_U.if_empty_n;
    assign fifo_intf_381.wr_en = AESL_inst_myproject.layer2_out_380_U.if_write & AESL_inst_myproject.layer2_out_380_U.if_full_n;
    assign fifo_intf_381.fifo_rd_block = 0;
    assign fifo_intf_381.fifo_wr_block = 0;
    assign fifo_intf_381.finish = finish;
    csv_file_dump fifo_csv_dumper_381;
    csv_file_dump cstatus_csv_dumper_381;
    df_fifo_monitor fifo_monitor_381;
    df_fifo_intf fifo_intf_382(clock,reset);
    assign fifo_intf_382.rd_en = AESL_inst_myproject.layer2_out_381_U.if_read & AESL_inst_myproject.layer2_out_381_U.if_empty_n;
    assign fifo_intf_382.wr_en = AESL_inst_myproject.layer2_out_381_U.if_write & AESL_inst_myproject.layer2_out_381_U.if_full_n;
    assign fifo_intf_382.fifo_rd_block = 0;
    assign fifo_intf_382.fifo_wr_block = 0;
    assign fifo_intf_382.finish = finish;
    csv_file_dump fifo_csv_dumper_382;
    csv_file_dump cstatus_csv_dumper_382;
    df_fifo_monitor fifo_monitor_382;
    df_fifo_intf fifo_intf_383(clock,reset);
    assign fifo_intf_383.rd_en = AESL_inst_myproject.layer2_out_382_U.if_read & AESL_inst_myproject.layer2_out_382_U.if_empty_n;
    assign fifo_intf_383.wr_en = AESL_inst_myproject.layer2_out_382_U.if_write & AESL_inst_myproject.layer2_out_382_U.if_full_n;
    assign fifo_intf_383.fifo_rd_block = 0;
    assign fifo_intf_383.fifo_wr_block = 0;
    assign fifo_intf_383.finish = finish;
    csv_file_dump fifo_csv_dumper_383;
    csv_file_dump cstatus_csv_dumper_383;
    df_fifo_monitor fifo_monitor_383;
    df_fifo_intf fifo_intf_384(clock,reset);
    assign fifo_intf_384.rd_en = AESL_inst_myproject.layer2_out_383_U.if_read & AESL_inst_myproject.layer2_out_383_U.if_empty_n;
    assign fifo_intf_384.wr_en = AESL_inst_myproject.layer2_out_383_U.if_write & AESL_inst_myproject.layer2_out_383_U.if_full_n;
    assign fifo_intf_384.fifo_rd_block = 0;
    assign fifo_intf_384.fifo_wr_block = 0;
    assign fifo_intf_384.finish = finish;
    csv_file_dump fifo_csv_dumper_384;
    csv_file_dump cstatus_csv_dumper_384;
    df_fifo_monitor fifo_monitor_384;
    df_fifo_intf fifo_intf_385(clock,reset);
    assign fifo_intf_385.rd_en = AESL_inst_myproject.layer2_out_384_U.if_read & AESL_inst_myproject.layer2_out_384_U.if_empty_n;
    assign fifo_intf_385.wr_en = AESL_inst_myproject.layer2_out_384_U.if_write & AESL_inst_myproject.layer2_out_384_U.if_full_n;
    assign fifo_intf_385.fifo_rd_block = 0;
    assign fifo_intf_385.fifo_wr_block = 0;
    assign fifo_intf_385.finish = finish;
    csv_file_dump fifo_csv_dumper_385;
    csv_file_dump cstatus_csv_dumper_385;
    df_fifo_monitor fifo_monitor_385;
    df_fifo_intf fifo_intf_386(clock,reset);
    assign fifo_intf_386.rd_en = AESL_inst_myproject.layer2_out_385_U.if_read & AESL_inst_myproject.layer2_out_385_U.if_empty_n;
    assign fifo_intf_386.wr_en = AESL_inst_myproject.layer2_out_385_U.if_write & AESL_inst_myproject.layer2_out_385_U.if_full_n;
    assign fifo_intf_386.fifo_rd_block = 0;
    assign fifo_intf_386.fifo_wr_block = 0;
    assign fifo_intf_386.finish = finish;
    csv_file_dump fifo_csv_dumper_386;
    csv_file_dump cstatus_csv_dumper_386;
    df_fifo_monitor fifo_monitor_386;
    df_fifo_intf fifo_intf_387(clock,reset);
    assign fifo_intf_387.rd_en = AESL_inst_myproject.layer2_out_386_U.if_read & AESL_inst_myproject.layer2_out_386_U.if_empty_n;
    assign fifo_intf_387.wr_en = AESL_inst_myproject.layer2_out_386_U.if_write & AESL_inst_myproject.layer2_out_386_U.if_full_n;
    assign fifo_intf_387.fifo_rd_block = 0;
    assign fifo_intf_387.fifo_wr_block = 0;
    assign fifo_intf_387.finish = finish;
    csv_file_dump fifo_csv_dumper_387;
    csv_file_dump cstatus_csv_dumper_387;
    df_fifo_monitor fifo_monitor_387;
    df_fifo_intf fifo_intf_388(clock,reset);
    assign fifo_intf_388.rd_en = AESL_inst_myproject.layer2_out_387_U.if_read & AESL_inst_myproject.layer2_out_387_U.if_empty_n;
    assign fifo_intf_388.wr_en = AESL_inst_myproject.layer2_out_387_U.if_write & AESL_inst_myproject.layer2_out_387_U.if_full_n;
    assign fifo_intf_388.fifo_rd_block = 0;
    assign fifo_intf_388.fifo_wr_block = 0;
    assign fifo_intf_388.finish = finish;
    csv_file_dump fifo_csv_dumper_388;
    csv_file_dump cstatus_csv_dumper_388;
    df_fifo_monitor fifo_monitor_388;
    df_fifo_intf fifo_intf_389(clock,reset);
    assign fifo_intf_389.rd_en = AESL_inst_myproject.layer2_out_388_U.if_read & AESL_inst_myproject.layer2_out_388_U.if_empty_n;
    assign fifo_intf_389.wr_en = AESL_inst_myproject.layer2_out_388_U.if_write & AESL_inst_myproject.layer2_out_388_U.if_full_n;
    assign fifo_intf_389.fifo_rd_block = 0;
    assign fifo_intf_389.fifo_wr_block = 0;
    assign fifo_intf_389.finish = finish;
    csv_file_dump fifo_csv_dumper_389;
    csv_file_dump cstatus_csv_dumper_389;
    df_fifo_monitor fifo_monitor_389;
    df_fifo_intf fifo_intf_390(clock,reset);
    assign fifo_intf_390.rd_en = AESL_inst_myproject.layer2_out_389_U.if_read & AESL_inst_myproject.layer2_out_389_U.if_empty_n;
    assign fifo_intf_390.wr_en = AESL_inst_myproject.layer2_out_389_U.if_write & AESL_inst_myproject.layer2_out_389_U.if_full_n;
    assign fifo_intf_390.fifo_rd_block = 0;
    assign fifo_intf_390.fifo_wr_block = 0;
    assign fifo_intf_390.finish = finish;
    csv_file_dump fifo_csv_dumper_390;
    csv_file_dump cstatus_csv_dumper_390;
    df_fifo_monitor fifo_monitor_390;
    df_fifo_intf fifo_intf_391(clock,reset);
    assign fifo_intf_391.rd_en = AESL_inst_myproject.layer2_out_390_U.if_read & AESL_inst_myproject.layer2_out_390_U.if_empty_n;
    assign fifo_intf_391.wr_en = AESL_inst_myproject.layer2_out_390_U.if_write & AESL_inst_myproject.layer2_out_390_U.if_full_n;
    assign fifo_intf_391.fifo_rd_block = 0;
    assign fifo_intf_391.fifo_wr_block = 0;
    assign fifo_intf_391.finish = finish;
    csv_file_dump fifo_csv_dumper_391;
    csv_file_dump cstatus_csv_dumper_391;
    df_fifo_monitor fifo_monitor_391;
    df_fifo_intf fifo_intf_392(clock,reset);
    assign fifo_intf_392.rd_en = AESL_inst_myproject.layer2_out_391_U.if_read & AESL_inst_myproject.layer2_out_391_U.if_empty_n;
    assign fifo_intf_392.wr_en = AESL_inst_myproject.layer2_out_391_U.if_write & AESL_inst_myproject.layer2_out_391_U.if_full_n;
    assign fifo_intf_392.fifo_rd_block = 0;
    assign fifo_intf_392.fifo_wr_block = 0;
    assign fifo_intf_392.finish = finish;
    csv_file_dump fifo_csv_dumper_392;
    csv_file_dump cstatus_csv_dumper_392;
    df_fifo_monitor fifo_monitor_392;
    df_fifo_intf fifo_intf_393(clock,reset);
    assign fifo_intf_393.rd_en = AESL_inst_myproject.layer2_out_392_U.if_read & AESL_inst_myproject.layer2_out_392_U.if_empty_n;
    assign fifo_intf_393.wr_en = AESL_inst_myproject.layer2_out_392_U.if_write & AESL_inst_myproject.layer2_out_392_U.if_full_n;
    assign fifo_intf_393.fifo_rd_block = 0;
    assign fifo_intf_393.fifo_wr_block = 0;
    assign fifo_intf_393.finish = finish;
    csv_file_dump fifo_csv_dumper_393;
    csv_file_dump cstatus_csv_dumper_393;
    df_fifo_monitor fifo_monitor_393;
    df_fifo_intf fifo_intf_394(clock,reset);
    assign fifo_intf_394.rd_en = AESL_inst_myproject.layer2_out_393_U.if_read & AESL_inst_myproject.layer2_out_393_U.if_empty_n;
    assign fifo_intf_394.wr_en = AESL_inst_myproject.layer2_out_393_U.if_write & AESL_inst_myproject.layer2_out_393_U.if_full_n;
    assign fifo_intf_394.fifo_rd_block = 0;
    assign fifo_intf_394.fifo_wr_block = 0;
    assign fifo_intf_394.finish = finish;
    csv_file_dump fifo_csv_dumper_394;
    csv_file_dump cstatus_csv_dumper_394;
    df_fifo_monitor fifo_monitor_394;
    df_fifo_intf fifo_intf_395(clock,reset);
    assign fifo_intf_395.rd_en = AESL_inst_myproject.layer2_out_394_U.if_read & AESL_inst_myproject.layer2_out_394_U.if_empty_n;
    assign fifo_intf_395.wr_en = AESL_inst_myproject.layer2_out_394_U.if_write & AESL_inst_myproject.layer2_out_394_U.if_full_n;
    assign fifo_intf_395.fifo_rd_block = 0;
    assign fifo_intf_395.fifo_wr_block = 0;
    assign fifo_intf_395.finish = finish;
    csv_file_dump fifo_csv_dumper_395;
    csv_file_dump cstatus_csv_dumper_395;
    df_fifo_monitor fifo_monitor_395;
    df_fifo_intf fifo_intf_396(clock,reset);
    assign fifo_intf_396.rd_en = AESL_inst_myproject.layer2_out_395_U.if_read & AESL_inst_myproject.layer2_out_395_U.if_empty_n;
    assign fifo_intf_396.wr_en = AESL_inst_myproject.layer2_out_395_U.if_write & AESL_inst_myproject.layer2_out_395_U.if_full_n;
    assign fifo_intf_396.fifo_rd_block = 0;
    assign fifo_intf_396.fifo_wr_block = 0;
    assign fifo_intf_396.finish = finish;
    csv_file_dump fifo_csv_dumper_396;
    csv_file_dump cstatus_csv_dumper_396;
    df_fifo_monitor fifo_monitor_396;
    df_fifo_intf fifo_intf_397(clock,reset);
    assign fifo_intf_397.rd_en = AESL_inst_myproject.layer2_out_396_U.if_read & AESL_inst_myproject.layer2_out_396_U.if_empty_n;
    assign fifo_intf_397.wr_en = AESL_inst_myproject.layer2_out_396_U.if_write & AESL_inst_myproject.layer2_out_396_U.if_full_n;
    assign fifo_intf_397.fifo_rd_block = 0;
    assign fifo_intf_397.fifo_wr_block = 0;
    assign fifo_intf_397.finish = finish;
    csv_file_dump fifo_csv_dumper_397;
    csv_file_dump cstatus_csv_dumper_397;
    df_fifo_monitor fifo_monitor_397;
    df_fifo_intf fifo_intf_398(clock,reset);
    assign fifo_intf_398.rd_en = AESL_inst_myproject.layer2_out_397_U.if_read & AESL_inst_myproject.layer2_out_397_U.if_empty_n;
    assign fifo_intf_398.wr_en = AESL_inst_myproject.layer2_out_397_U.if_write & AESL_inst_myproject.layer2_out_397_U.if_full_n;
    assign fifo_intf_398.fifo_rd_block = 0;
    assign fifo_intf_398.fifo_wr_block = 0;
    assign fifo_intf_398.finish = finish;
    csv_file_dump fifo_csv_dumper_398;
    csv_file_dump cstatus_csv_dumper_398;
    df_fifo_monitor fifo_monitor_398;
    df_fifo_intf fifo_intf_399(clock,reset);
    assign fifo_intf_399.rd_en = AESL_inst_myproject.layer2_out_398_U.if_read & AESL_inst_myproject.layer2_out_398_U.if_empty_n;
    assign fifo_intf_399.wr_en = AESL_inst_myproject.layer2_out_398_U.if_write & AESL_inst_myproject.layer2_out_398_U.if_full_n;
    assign fifo_intf_399.fifo_rd_block = 0;
    assign fifo_intf_399.fifo_wr_block = 0;
    assign fifo_intf_399.finish = finish;
    csv_file_dump fifo_csv_dumper_399;
    csv_file_dump cstatus_csv_dumper_399;
    df_fifo_monitor fifo_monitor_399;
    df_fifo_intf fifo_intf_400(clock,reset);
    assign fifo_intf_400.rd_en = AESL_inst_myproject.layer2_out_399_U.if_read & AESL_inst_myproject.layer2_out_399_U.if_empty_n;
    assign fifo_intf_400.wr_en = AESL_inst_myproject.layer2_out_399_U.if_write & AESL_inst_myproject.layer2_out_399_U.if_full_n;
    assign fifo_intf_400.fifo_rd_block = 0;
    assign fifo_intf_400.fifo_wr_block = 0;
    assign fifo_intf_400.finish = finish;
    csv_file_dump fifo_csv_dumper_400;
    csv_file_dump cstatus_csv_dumper_400;
    df_fifo_monitor fifo_monitor_400;
    df_fifo_intf fifo_intf_401(clock,reset);
    assign fifo_intf_401.rd_en = AESL_inst_myproject.layer2_out_400_U.if_read & AESL_inst_myproject.layer2_out_400_U.if_empty_n;
    assign fifo_intf_401.wr_en = AESL_inst_myproject.layer2_out_400_U.if_write & AESL_inst_myproject.layer2_out_400_U.if_full_n;
    assign fifo_intf_401.fifo_rd_block = 0;
    assign fifo_intf_401.fifo_wr_block = 0;
    assign fifo_intf_401.finish = finish;
    csv_file_dump fifo_csv_dumper_401;
    csv_file_dump cstatus_csv_dumper_401;
    df_fifo_monitor fifo_monitor_401;
    df_fifo_intf fifo_intf_402(clock,reset);
    assign fifo_intf_402.rd_en = AESL_inst_myproject.layer2_out_401_U.if_read & AESL_inst_myproject.layer2_out_401_U.if_empty_n;
    assign fifo_intf_402.wr_en = AESL_inst_myproject.layer2_out_401_U.if_write & AESL_inst_myproject.layer2_out_401_U.if_full_n;
    assign fifo_intf_402.fifo_rd_block = 0;
    assign fifo_intf_402.fifo_wr_block = 0;
    assign fifo_intf_402.finish = finish;
    csv_file_dump fifo_csv_dumper_402;
    csv_file_dump cstatus_csv_dumper_402;
    df_fifo_monitor fifo_monitor_402;
    df_fifo_intf fifo_intf_403(clock,reset);
    assign fifo_intf_403.rd_en = AESL_inst_myproject.layer2_out_402_U.if_read & AESL_inst_myproject.layer2_out_402_U.if_empty_n;
    assign fifo_intf_403.wr_en = AESL_inst_myproject.layer2_out_402_U.if_write & AESL_inst_myproject.layer2_out_402_U.if_full_n;
    assign fifo_intf_403.fifo_rd_block = 0;
    assign fifo_intf_403.fifo_wr_block = 0;
    assign fifo_intf_403.finish = finish;
    csv_file_dump fifo_csv_dumper_403;
    csv_file_dump cstatus_csv_dumper_403;
    df_fifo_monitor fifo_monitor_403;
    df_fifo_intf fifo_intf_404(clock,reset);
    assign fifo_intf_404.rd_en = AESL_inst_myproject.layer2_out_403_U.if_read & AESL_inst_myproject.layer2_out_403_U.if_empty_n;
    assign fifo_intf_404.wr_en = AESL_inst_myproject.layer2_out_403_U.if_write & AESL_inst_myproject.layer2_out_403_U.if_full_n;
    assign fifo_intf_404.fifo_rd_block = 0;
    assign fifo_intf_404.fifo_wr_block = 0;
    assign fifo_intf_404.finish = finish;
    csv_file_dump fifo_csv_dumper_404;
    csv_file_dump cstatus_csv_dumper_404;
    df_fifo_monitor fifo_monitor_404;
    df_fifo_intf fifo_intf_405(clock,reset);
    assign fifo_intf_405.rd_en = AESL_inst_myproject.layer2_out_404_U.if_read & AESL_inst_myproject.layer2_out_404_U.if_empty_n;
    assign fifo_intf_405.wr_en = AESL_inst_myproject.layer2_out_404_U.if_write & AESL_inst_myproject.layer2_out_404_U.if_full_n;
    assign fifo_intf_405.fifo_rd_block = 0;
    assign fifo_intf_405.fifo_wr_block = 0;
    assign fifo_intf_405.finish = finish;
    csv_file_dump fifo_csv_dumper_405;
    csv_file_dump cstatus_csv_dumper_405;
    df_fifo_monitor fifo_monitor_405;
    df_fifo_intf fifo_intf_406(clock,reset);
    assign fifo_intf_406.rd_en = AESL_inst_myproject.layer2_out_405_U.if_read & AESL_inst_myproject.layer2_out_405_U.if_empty_n;
    assign fifo_intf_406.wr_en = AESL_inst_myproject.layer2_out_405_U.if_write & AESL_inst_myproject.layer2_out_405_U.if_full_n;
    assign fifo_intf_406.fifo_rd_block = 0;
    assign fifo_intf_406.fifo_wr_block = 0;
    assign fifo_intf_406.finish = finish;
    csv_file_dump fifo_csv_dumper_406;
    csv_file_dump cstatus_csv_dumper_406;
    df_fifo_monitor fifo_monitor_406;
    df_fifo_intf fifo_intf_407(clock,reset);
    assign fifo_intf_407.rd_en = AESL_inst_myproject.layer2_out_406_U.if_read & AESL_inst_myproject.layer2_out_406_U.if_empty_n;
    assign fifo_intf_407.wr_en = AESL_inst_myproject.layer2_out_406_U.if_write & AESL_inst_myproject.layer2_out_406_U.if_full_n;
    assign fifo_intf_407.fifo_rd_block = 0;
    assign fifo_intf_407.fifo_wr_block = 0;
    assign fifo_intf_407.finish = finish;
    csv_file_dump fifo_csv_dumper_407;
    csv_file_dump cstatus_csv_dumper_407;
    df_fifo_monitor fifo_monitor_407;
    df_fifo_intf fifo_intf_408(clock,reset);
    assign fifo_intf_408.rd_en = AESL_inst_myproject.layer2_out_407_U.if_read & AESL_inst_myproject.layer2_out_407_U.if_empty_n;
    assign fifo_intf_408.wr_en = AESL_inst_myproject.layer2_out_407_U.if_write & AESL_inst_myproject.layer2_out_407_U.if_full_n;
    assign fifo_intf_408.fifo_rd_block = 0;
    assign fifo_intf_408.fifo_wr_block = 0;
    assign fifo_intf_408.finish = finish;
    csv_file_dump fifo_csv_dumper_408;
    csv_file_dump cstatus_csv_dumper_408;
    df_fifo_monitor fifo_monitor_408;
    df_fifo_intf fifo_intf_409(clock,reset);
    assign fifo_intf_409.rd_en = AESL_inst_myproject.layer2_out_408_U.if_read & AESL_inst_myproject.layer2_out_408_U.if_empty_n;
    assign fifo_intf_409.wr_en = AESL_inst_myproject.layer2_out_408_U.if_write & AESL_inst_myproject.layer2_out_408_U.if_full_n;
    assign fifo_intf_409.fifo_rd_block = 0;
    assign fifo_intf_409.fifo_wr_block = 0;
    assign fifo_intf_409.finish = finish;
    csv_file_dump fifo_csv_dumper_409;
    csv_file_dump cstatus_csv_dumper_409;
    df_fifo_monitor fifo_monitor_409;
    df_fifo_intf fifo_intf_410(clock,reset);
    assign fifo_intf_410.rd_en = AESL_inst_myproject.layer2_out_409_U.if_read & AESL_inst_myproject.layer2_out_409_U.if_empty_n;
    assign fifo_intf_410.wr_en = AESL_inst_myproject.layer2_out_409_U.if_write & AESL_inst_myproject.layer2_out_409_U.if_full_n;
    assign fifo_intf_410.fifo_rd_block = 0;
    assign fifo_intf_410.fifo_wr_block = 0;
    assign fifo_intf_410.finish = finish;
    csv_file_dump fifo_csv_dumper_410;
    csv_file_dump cstatus_csv_dumper_410;
    df_fifo_monitor fifo_monitor_410;
    df_fifo_intf fifo_intf_411(clock,reset);
    assign fifo_intf_411.rd_en = AESL_inst_myproject.layer2_out_410_U.if_read & AESL_inst_myproject.layer2_out_410_U.if_empty_n;
    assign fifo_intf_411.wr_en = AESL_inst_myproject.layer2_out_410_U.if_write & AESL_inst_myproject.layer2_out_410_U.if_full_n;
    assign fifo_intf_411.fifo_rd_block = 0;
    assign fifo_intf_411.fifo_wr_block = 0;
    assign fifo_intf_411.finish = finish;
    csv_file_dump fifo_csv_dumper_411;
    csv_file_dump cstatus_csv_dumper_411;
    df_fifo_monitor fifo_monitor_411;
    df_fifo_intf fifo_intf_412(clock,reset);
    assign fifo_intf_412.rd_en = AESL_inst_myproject.layer2_out_411_U.if_read & AESL_inst_myproject.layer2_out_411_U.if_empty_n;
    assign fifo_intf_412.wr_en = AESL_inst_myproject.layer2_out_411_U.if_write & AESL_inst_myproject.layer2_out_411_U.if_full_n;
    assign fifo_intf_412.fifo_rd_block = 0;
    assign fifo_intf_412.fifo_wr_block = 0;
    assign fifo_intf_412.finish = finish;
    csv_file_dump fifo_csv_dumper_412;
    csv_file_dump cstatus_csv_dumper_412;
    df_fifo_monitor fifo_monitor_412;
    df_fifo_intf fifo_intf_413(clock,reset);
    assign fifo_intf_413.rd_en = AESL_inst_myproject.layer2_out_412_U.if_read & AESL_inst_myproject.layer2_out_412_U.if_empty_n;
    assign fifo_intf_413.wr_en = AESL_inst_myproject.layer2_out_412_U.if_write & AESL_inst_myproject.layer2_out_412_U.if_full_n;
    assign fifo_intf_413.fifo_rd_block = 0;
    assign fifo_intf_413.fifo_wr_block = 0;
    assign fifo_intf_413.finish = finish;
    csv_file_dump fifo_csv_dumper_413;
    csv_file_dump cstatus_csv_dumper_413;
    df_fifo_monitor fifo_monitor_413;
    df_fifo_intf fifo_intf_414(clock,reset);
    assign fifo_intf_414.rd_en = AESL_inst_myproject.layer2_out_413_U.if_read & AESL_inst_myproject.layer2_out_413_U.if_empty_n;
    assign fifo_intf_414.wr_en = AESL_inst_myproject.layer2_out_413_U.if_write & AESL_inst_myproject.layer2_out_413_U.if_full_n;
    assign fifo_intf_414.fifo_rd_block = 0;
    assign fifo_intf_414.fifo_wr_block = 0;
    assign fifo_intf_414.finish = finish;
    csv_file_dump fifo_csv_dumper_414;
    csv_file_dump cstatus_csv_dumper_414;
    df_fifo_monitor fifo_monitor_414;
    df_fifo_intf fifo_intf_415(clock,reset);
    assign fifo_intf_415.rd_en = AESL_inst_myproject.layer2_out_414_U.if_read & AESL_inst_myproject.layer2_out_414_U.if_empty_n;
    assign fifo_intf_415.wr_en = AESL_inst_myproject.layer2_out_414_U.if_write & AESL_inst_myproject.layer2_out_414_U.if_full_n;
    assign fifo_intf_415.fifo_rd_block = 0;
    assign fifo_intf_415.fifo_wr_block = 0;
    assign fifo_intf_415.finish = finish;
    csv_file_dump fifo_csv_dumper_415;
    csv_file_dump cstatus_csv_dumper_415;
    df_fifo_monitor fifo_monitor_415;
    df_fifo_intf fifo_intf_416(clock,reset);
    assign fifo_intf_416.rd_en = AESL_inst_myproject.layer2_out_415_U.if_read & AESL_inst_myproject.layer2_out_415_U.if_empty_n;
    assign fifo_intf_416.wr_en = AESL_inst_myproject.layer2_out_415_U.if_write & AESL_inst_myproject.layer2_out_415_U.if_full_n;
    assign fifo_intf_416.fifo_rd_block = 0;
    assign fifo_intf_416.fifo_wr_block = 0;
    assign fifo_intf_416.finish = finish;
    csv_file_dump fifo_csv_dumper_416;
    csv_file_dump cstatus_csv_dumper_416;
    df_fifo_monitor fifo_monitor_416;
    df_fifo_intf fifo_intf_417(clock,reset);
    assign fifo_intf_417.rd_en = AESL_inst_myproject.layer2_out_416_U.if_read & AESL_inst_myproject.layer2_out_416_U.if_empty_n;
    assign fifo_intf_417.wr_en = AESL_inst_myproject.layer2_out_416_U.if_write & AESL_inst_myproject.layer2_out_416_U.if_full_n;
    assign fifo_intf_417.fifo_rd_block = 0;
    assign fifo_intf_417.fifo_wr_block = 0;
    assign fifo_intf_417.finish = finish;
    csv_file_dump fifo_csv_dumper_417;
    csv_file_dump cstatus_csv_dumper_417;
    df_fifo_monitor fifo_monitor_417;
    df_fifo_intf fifo_intf_418(clock,reset);
    assign fifo_intf_418.rd_en = AESL_inst_myproject.layer2_out_417_U.if_read & AESL_inst_myproject.layer2_out_417_U.if_empty_n;
    assign fifo_intf_418.wr_en = AESL_inst_myproject.layer2_out_417_U.if_write & AESL_inst_myproject.layer2_out_417_U.if_full_n;
    assign fifo_intf_418.fifo_rd_block = 0;
    assign fifo_intf_418.fifo_wr_block = 0;
    assign fifo_intf_418.finish = finish;
    csv_file_dump fifo_csv_dumper_418;
    csv_file_dump cstatus_csv_dumper_418;
    df_fifo_monitor fifo_monitor_418;
    df_fifo_intf fifo_intf_419(clock,reset);
    assign fifo_intf_419.rd_en = AESL_inst_myproject.layer2_out_418_U.if_read & AESL_inst_myproject.layer2_out_418_U.if_empty_n;
    assign fifo_intf_419.wr_en = AESL_inst_myproject.layer2_out_418_U.if_write & AESL_inst_myproject.layer2_out_418_U.if_full_n;
    assign fifo_intf_419.fifo_rd_block = 0;
    assign fifo_intf_419.fifo_wr_block = 0;
    assign fifo_intf_419.finish = finish;
    csv_file_dump fifo_csv_dumper_419;
    csv_file_dump cstatus_csv_dumper_419;
    df_fifo_monitor fifo_monitor_419;
    df_fifo_intf fifo_intf_420(clock,reset);
    assign fifo_intf_420.rd_en = AESL_inst_myproject.layer2_out_419_U.if_read & AESL_inst_myproject.layer2_out_419_U.if_empty_n;
    assign fifo_intf_420.wr_en = AESL_inst_myproject.layer2_out_419_U.if_write & AESL_inst_myproject.layer2_out_419_U.if_full_n;
    assign fifo_intf_420.fifo_rd_block = 0;
    assign fifo_intf_420.fifo_wr_block = 0;
    assign fifo_intf_420.finish = finish;
    csv_file_dump fifo_csv_dumper_420;
    csv_file_dump cstatus_csv_dumper_420;
    df_fifo_monitor fifo_monitor_420;
    df_fifo_intf fifo_intf_421(clock,reset);
    assign fifo_intf_421.rd_en = AESL_inst_myproject.layer2_out_420_U.if_read & AESL_inst_myproject.layer2_out_420_U.if_empty_n;
    assign fifo_intf_421.wr_en = AESL_inst_myproject.layer2_out_420_U.if_write & AESL_inst_myproject.layer2_out_420_U.if_full_n;
    assign fifo_intf_421.fifo_rd_block = 0;
    assign fifo_intf_421.fifo_wr_block = 0;
    assign fifo_intf_421.finish = finish;
    csv_file_dump fifo_csv_dumper_421;
    csv_file_dump cstatus_csv_dumper_421;
    df_fifo_monitor fifo_monitor_421;
    df_fifo_intf fifo_intf_422(clock,reset);
    assign fifo_intf_422.rd_en = AESL_inst_myproject.layer2_out_421_U.if_read & AESL_inst_myproject.layer2_out_421_U.if_empty_n;
    assign fifo_intf_422.wr_en = AESL_inst_myproject.layer2_out_421_U.if_write & AESL_inst_myproject.layer2_out_421_U.if_full_n;
    assign fifo_intf_422.fifo_rd_block = 0;
    assign fifo_intf_422.fifo_wr_block = 0;
    assign fifo_intf_422.finish = finish;
    csv_file_dump fifo_csv_dumper_422;
    csv_file_dump cstatus_csv_dumper_422;
    df_fifo_monitor fifo_monitor_422;
    df_fifo_intf fifo_intf_423(clock,reset);
    assign fifo_intf_423.rd_en = AESL_inst_myproject.layer2_out_422_U.if_read & AESL_inst_myproject.layer2_out_422_U.if_empty_n;
    assign fifo_intf_423.wr_en = AESL_inst_myproject.layer2_out_422_U.if_write & AESL_inst_myproject.layer2_out_422_U.if_full_n;
    assign fifo_intf_423.fifo_rd_block = 0;
    assign fifo_intf_423.fifo_wr_block = 0;
    assign fifo_intf_423.finish = finish;
    csv_file_dump fifo_csv_dumper_423;
    csv_file_dump cstatus_csv_dumper_423;
    df_fifo_monitor fifo_monitor_423;
    df_fifo_intf fifo_intf_424(clock,reset);
    assign fifo_intf_424.rd_en = AESL_inst_myproject.layer2_out_423_U.if_read & AESL_inst_myproject.layer2_out_423_U.if_empty_n;
    assign fifo_intf_424.wr_en = AESL_inst_myproject.layer2_out_423_U.if_write & AESL_inst_myproject.layer2_out_423_U.if_full_n;
    assign fifo_intf_424.fifo_rd_block = 0;
    assign fifo_intf_424.fifo_wr_block = 0;
    assign fifo_intf_424.finish = finish;
    csv_file_dump fifo_csv_dumper_424;
    csv_file_dump cstatus_csv_dumper_424;
    df_fifo_monitor fifo_monitor_424;
    df_fifo_intf fifo_intf_425(clock,reset);
    assign fifo_intf_425.rd_en = AESL_inst_myproject.layer2_out_424_U.if_read & AESL_inst_myproject.layer2_out_424_U.if_empty_n;
    assign fifo_intf_425.wr_en = AESL_inst_myproject.layer2_out_424_U.if_write & AESL_inst_myproject.layer2_out_424_U.if_full_n;
    assign fifo_intf_425.fifo_rd_block = 0;
    assign fifo_intf_425.fifo_wr_block = 0;
    assign fifo_intf_425.finish = finish;
    csv_file_dump fifo_csv_dumper_425;
    csv_file_dump cstatus_csv_dumper_425;
    df_fifo_monitor fifo_monitor_425;
    df_fifo_intf fifo_intf_426(clock,reset);
    assign fifo_intf_426.rd_en = AESL_inst_myproject.layer2_out_425_U.if_read & AESL_inst_myproject.layer2_out_425_U.if_empty_n;
    assign fifo_intf_426.wr_en = AESL_inst_myproject.layer2_out_425_U.if_write & AESL_inst_myproject.layer2_out_425_U.if_full_n;
    assign fifo_intf_426.fifo_rd_block = 0;
    assign fifo_intf_426.fifo_wr_block = 0;
    assign fifo_intf_426.finish = finish;
    csv_file_dump fifo_csv_dumper_426;
    csv_file_dump cstatus_csv_dumper_426;
    df_fifo_monitor fifo_monitor_426;
    df_fifo_intf fifo_intf_427(clock,reset);
    assign fifo_intf_427.rd_en = AESL_inst_myproject.layer2_out_426_U.if_read & AESL_inst_myproject.layer2_out_426_U.if_empty_n;
    assign fifo_intf_427.wr_en = AESL_inst_myproject.layer2_out_426_U.if_write & AESL_inst_myproject.layer2_out_426_U.if_full_n;
    assign fifo_intf_427.fifo_rd_block = 0;
    assign fifo_intf_427.fifo_wr_block = 0;
    assign fifo_intf_427.finish = finish;
    csv_file_dump fifo_csv_dumper_427;
    csv_file_dump cstatus_csv_dumper_427;
    df_fifo_monitor fifo_monitor_427;
    df_fifo_intf fifo_intf_428(clock,reset);
    assign fifo_intf_428.rd_en = AESL_inst_myproject.layer2_out_427_U.if_read & AESL_inst_myproject.layer2_out_427_U.if_empty_n;
    assign fifo_intf_428.wr_en = AESL_inst_myproject.layer2_out_427_U.if_write & AESL_inst_myproject.layer2_out_427_U.if_full_n;
    assign fifo_intf_428.fifo_rd_block = 0;
    assign fifo_intf_428.fifo_wr_block = 0;
    assign fifo_intf_428.finish = finish;
    csv_file_dump fifo_csv_dumper_428;
    csv_file_dump cstatus_csv_dumper_428;
    df_fifo_monitor fifo_monitor_428;
    df_fifo_intf fifo_intf_429(clock,reset);
    assign fifo_intf_429.rd_en = AESL_inst_myproject.layer2_out_428_U.if_read & AESL_inst_myproject.layer2_out_428_U.if_empty_n;
    assign fifo_intf_429.wr_en = AESL_inst_myproject.layer2_out_428_U.if_write & AESL_inst_myproject.layer2_out_428_U.if_full_n;
    assign fifo_intf_429.fifo_rd_block = 0;
    assign fifo_intf_429.fifo_wr_block = 0;
    assign fifo_intf_429.finish = finish;
    csv_file_dump fifo_csv_dumper_429;
    csv_file_dump cstatus_csv_dumper_429;
    df_fifo_monitor fifo_monitor_429;
    df_fifo_intf fifo_intf_430(clock,reset);
    assign fifo_intf_430.rd_en = AESL_inst_myproject.layer2_out_429_U.if_read & AESL_inst_myproject.layer2_out_429_U.if_empty_n;
    assign fifo_intf_430.wr_en = AESL_inst_myproject.layer2_out_429_U.if_write & AESL_inst_myproject.layer2_out_429_U.if_full_n;
    assign fifo_intf_430.fifo_rd_block = 0;
    assign fifo_intf_430.fifo_wr_block = 0;
    assign fifo_intf_430.finish = finish;
    csv_file_dump fifo_csv_dumper_430;
    csv_file_dump cstatus_csv_dumper_430;
    df_fifo_monitor fifo_monitor_430;
    df_fifo_intf fifo_intf_431(clock,reset);
    assign fifo_intf_431.rd_en = AESL_inst_myproject.layer2_out_430_U.if_read & AESL_inst_myproject.layer2_out_430_U.if_empty_n;
    assign fifo_intf_431.wr_en = AESL_inst_myproject.layer2_out_430_U.if_write & AESL_inst_myproject.layer2_out_430_U.if_full_n;
    assign fifo_intf_431.fifo_rd_block = 0;
    assign fifo_intf_431.fifo_wr_block = 0;
    assign fifo_intf_431.finish = finish;
    csv_file_dump fifo_csv_dumper_431;
    csv_file_dump cstatus_csv_dumper_431;
    df_fifo_monitor fifo_monitor_431;
    df_fifo_intf fifo_intf_432(clock,reset);
    assign fifo_intf_432.rd_en = AESL_inst_myproject.layer2_out_431_U.if_read & AESL_inst_myproject.layer2_out_431_U.if_empty_n;
    assign fifo_intf_432.wr_en = AESL_inst_myproject.layer2_out_431_U.if_write & AESL_inst_myproject.layer2_out_431_U.if_full_n;
    assign fifo_intf_432.fifo_rd_block = 0;
    assign fifo_intf_432.fifo_wr_block = 0;
    assign fifo_intf_432.finish = finish;
    csv_file_dump fifo_csv_dumper_432;
    csv_file_dump cstatus_csv_dumper_432;
    df_fifo_monitor fifo_monitor_432;
    df_fifo_intf fifo_intf_433(clock,reset);
    assign fifo_intf_433.rd_en = AESL_inst_myproject.layer2_out_432_U.if_read & AESL_inst_myproject.layer2_out_432_U.if_empty_n;
    assign fifo_intf_433.wr_en = AESL_inst_myproject.layer2_out_432_U.if_write & AESL_inst_myproject.layer2_out_432_U.if_full_n;
    assign fifo_intf_433.fifo_rd_block = 0;
    assign fifo_intf_433.fifo_wr_block = 0;
    assign fifo_intf_433.finish = finish;
    csv_file_dump fifo_csv_dumper_433;
    csv_file_dump cstatus_csv_dumper_433;
    df_fifo_monitor fifo_monitor_433;
    df_fifo_intf fifo_intf_434(clock,reset);
    assign fifo_intf_434.rd_en = AESL_inst_myproject.layer2_out_433_U.if_read & AESL_inst_myproject.layer2_out_433_U.if_empty_n;
    assign fifo_intf_434.wr_en = AESL_inst_myproject.layer2_out_433_U.if_write & AESL_inst_myproject.layer2_out_433_U.if_full_n;
    assign fifo_intf_434.fifo_rd_block = 0;
    assign fifo_intf_434.fifo_wr_block = 0;
    assign fifo_intf_434.finish = finish;
    csv_file_dump fifo_csv_dumper_434;
    csv_file_dump cstatus_csv_dumper_434;
    df_fifo_monitor fifo_monitor_434;
    df_fifo_intf fifo_intf_435(clock,reset);
    assign fifo_intf_435.rd_en = AESL_inst_myproject.layer2_out_434_U.if_read & AESL_inst_myproject.layer2_out_434_U.if_empty_n;
    assign fifo_intf_435.wr_en = AESL_inst_myproject.layer2_out_434_U.if_write & AESL_inst_myproject.layer2_out_434_U.if_full_n;
    assign fifo_intf_435.fifo_rd_block = 0;
    assign fifo_intf_435.fifo_wr_block = 0;
    assign fifo_intf_435.finish = finish;
    csv_file_dump fifo_csv_dumper_435;
    csv_file_dump cstatus_csv_dumper_435;
    df_fifo_monitor fifo_monitor_435;
    df_fifo_intf fifo_intf_436(clock,reset);
    assign fifo_intf_436.rd_en = AESL_inst_myproject.layer2_out_435_U.if_read & AESL_inst_myproject.layer2_out_435_U.if_empty_n;
    assign fifo_intf_436.wr_en = AESL_inst_myproject.layer2_out_435_U.if_write & AESL_inst_myproject.layer2_out_435_U.if_full_n;
    assign fifo_intf_436.fifo_rd_block = 0;
    assign fifo_intf_436.fifo_wr_block = 0;
    assign fifo_intf_436.finish = finish;
    csv_file_dump fifo_csv_dumper_436;
    csv_file_dump cstatus_csv_dumper_436;
    df_fifo_monitor fifo_monitor_436;
    df_fifo_intf fifo_intf_437(clock,reset);
    assign fifo_intf_437.rd_en = AESL_inst_myproject.layer2_out_436_U.if_read & AESL_inst_myproject.layer2_out_436_U.if_empty_n;
    assign fifo_intf_437.wr_en = AESL_inst_myproject.layer2_out_436_U.if_write & AESL_inst_myproject.layer2_out_436_U.if_full_n;
    assign fifo_intf_437.fifo_rd_block = 0;
    assign fifo_intf_437.fifo_wr_block = 0;
    assign fifo_intf_437.finish = finish;
    csv_file_dump fifo_csv_dumper_437;
    csv_file_dump cstatus_csv_dumper_437;
    df_fifo_monitor fifo_monitor_437;
    df_fifo_intf fifo_intf_438(clock,reset);
    assign fifo_intf_438.rd_en = AESL_inst_myproject.layer2_out_437_U.if_read & AESL_inst_myproject.layer2_out_437_U.if_empty_n;
    assign fifo_intf_438.wr_en = AESL_inst_myproject.layer2_out_437_U.if_write & AESL_inst_myproject.layer2_out_437_U.if_full_n;
    assign fifo_intf_438.fifo_rd_block = 0;
    assign fifo_intf_438.fifo_wr_block = 0;
    assign fifo_intf_438.finish = finish;
    csv_file_dump fifo_csv_dumper_438;
    csv_file_dump cstatus_csv_dumper_438;
    df_fifo_monitor fifo_monitor_438;
    df_fifo_intf fifo_intf_439(clock,reset);
    assign fifo_intf_439.rd_en = AESL_inst_myproject.layer2_out_438_U.if_read & AESL_inst_myproject.layer2_out_438_U.if_empty_n;
    assign fifo_intf_439.wr_en = AESL_inst_myproject.layer2_out_438_U.if_write & AESL_inst_myproject.layer2_out_438_U.if_full_n;
    assign fifo_intf_439.fifo_rd_block = 0;
    assign fifo_intf_439.fifo_wr_block = 0;
    assign fifo_intf_439.finish = finish;
    csv_file_dump fifo_csv_dumper_439;
    csv_file_dump cstatus_csv_dumper_439;
    df_fifo_monitor fifo_monitor_439;
    df_fifo_intf fifo_intf_440(clock,reset);
    assign fifo_intf_440.rd_en = AESL_inst_myproject.layer2_out_439_U.if_read & AESL_inst_myproject.layer2_out_439_U.if_empty_n;
    assign fifo_intf_440.wr_en = AESL_inst_myproject.layer2_out_439_U.if_write & AESL_inst_myproject.layer2_out_439_U.if_full_n;
    assign fifo_intf_440.fifo_rd_block = 0;
    assign fifo_intf_440.fifo_wr_block = 0;
    assign fifo_intf_440.finish = finish;
    csv_file_dump fifo_csv_dumper_440;
    csv_file_dump cstatus_csv_dumper_440;
    df_fifo_monitor fifo_monitor_440;
    df_fifo_intf fifo_intf_441(clock,reset);
    assign fifo_intf_441.rd_en = AESL_inst_myproject.layer2_out_440_U.if_read & AESL_inst_myproject.layer2_out_440_U.if_empty_n;
    assign fifo_intf_441.wr_en = AESL_inst_myproject.layer2_out_440_U.if_write & AESL_inst_myproject.layer2_out_440_U.if_full_n;
    assign fifo_intf_441.fifo_rd_block = 0;
    assign fifo_intf_441.fifo_wr_block = 0;
    assign fifo_intf_441.finish = finish;
    csv_file_dump fifo_csv_dumper_441;
    csv_file_dump cstatus_csv_dumper_441;
    df_fifo_monitor fifo_monitor_441;
    df_fifo_intf fifo_intf_442(clock,reset);
    assign fifo_intf_442.rd_en = AESL_inst_myproject.layer2_out_441_U.if_read & AESL_inst_myproject.layer2_out_441_U.if_empty_n;
    assign fifo_intf_442.wr_en = AESL_inst_myproject.layer2_out_441_U.if_write & AESL_inst_myproject.layer2_out_441_U.if_full_n;
    assign fifo_intf_442.fifo_rd_block = 0;
    assign fifo_intf_442.fifo_wr_block = 0;
    assign fifo_intf_442.finish = finish;
    csv_file_dump fifo_csv_dumper_442;
    csv_file_dump cstatus_csv_dumper_442;
    df_fifo_monitor fifo_monitor_442;
    df_fifo_intf fifo_intf_443(clock,reset);
    assign fifo_intf_443.rd_en = AESL_inst_myproject.layer2_out_442_U.if_read & AESL_inst_myproject.layer2_out_442_U.if_empty_n;
    assign fifo_intf_443.wr_en = AESL_inst_myproject.layer2_out_442_U.if_write & AESL_inst_myproject.layer2_out_442_U.if_full_n;
    assign fifo_intf_443.fifo_rd_block = 0;
    assign fifo_intf_443.fifo_wr_block = 0;
    assign fifo_intf_443.finish = finish;
    csv_file_dump fifo_csv_dumper_443;
    csv_file_dump cstatus_csv_dumper_443;
    df_fifo_monitor fifo_monitor_443;
    df_fifo_intf fifo_intf_444(clock,reset);
    assign fifo_intf_444.rd_en = AESL_inst_myproject.layer2_out_443_U.if_read & AESL_inst_myproject.layer2_out_443_U.if_empty_n;
    assign fifo_intf_444.wr_en = AESL_inst_myproject.layer2_out_443_U.if_write & AESL_inst_myproject.layer2_out_443_U.if_full_n;
    assign fifo_intf_444.fifo_rd_block = 0;
    assign fifo_intf_444.fifo_wr_block = 0;
    assign fifo_intf_444.finish = finish;
    csv_file_dump fifo_csv_dumper_444;
    csv_file_dump cstatus_csv_dumper_444;
    df_fifo_monitor fifo_monitor_444;
    df_fifo_intf fifo_intf_445(clock,reset);
    assign fifo_intf_445.rd_en = AESL_inst_myproject.layer2_out_444_U.if_read & AESL_inst_myproject.layer2_out_444_U.if_empty_n;
    assign fifo_intf_445.wr_en = AESL_inst_myproject.layer2_out_444_U.if_write & AESL_inst_myproject.layer2_out_444_U.if_full_n;
    assign fifo_intf_445.fifo_rd_block = 0;
    assign fifo_intf_445.fifo_wr_block = 0;
    assign fifo_intf_445.finish = finish;
    csv_file_dump fifo_csv_dumper_445;
    csv_file_dump cstatus_csv_dumper_445;
    df_fifo_monitor fifo_monitor_445;
    df_fifo_intf fifo_intf_446(clock,reset);
    assign fifo_intf_446.rd_en = AESL_inst_myproject.layer2_out_445_U.if_read & AESL_inst_myproject.layer2_out_445_U.if_empty_n;
    assign fifo_intf_446.wr_en = AESL_inst_myproject.layer2_out_445_U.if_write & AESL_inst_myproject.layer2_out_445_U.if_full_n;
    assign fifo_intf_446.fifo_rd_block = 0;
    assign fifo_intf_446.fifo_wr_block = 0;
    assign fifo_intf_446.finish = finish;
    csv_file_dump fifo_csv_dumper_446;
    csv_file_dump cstatus_csv_dumper_446;
    df_fifo_monitor fifo_monitor_446;
    df_fifo_intf fifo_intf_447(clock,reset);
    assign fifo_intf_447.rd_en = AESL_inst_myproject.layer2_out_446_U.if_read & AESL_inst_myproject.layer2_out_446_U.if_empty_n;
    assign fifo_intf_447.wr_en = AESL_inst_myproject.layer2_out_446_U.if_write & AESL_inst_myproject.layer2_out_446_U.if_full_n;
    assign fifo_intf_447.fifo_rd_block = 0;
    assign fifo_intf_447.fifo_wr_block = 0;
    assign fifo_intf_447.finish = finish;
    csv_file_dump fifo_csv_dumper_447;
    csv_file_dump cstatus_csv_dumper_447;
    df_fifo_monitor fifo_monitor_447;
    df_fifo_intf fifo_intf_448(clock,reset);
    assign fifo_intf_448.rd_en = AESL_inst_myproject.layer2_out_447_U.if_read & AESL_inst_myproject.layer2_out_447_U.if_empty_n;
    assign fifo_intf_448.wr_en = AESL_inst_myproject.layer2_out_447_U.if_write & AESL_inst_myproject.layer2_out_447_U.if_full_n;
    assign fifo_intf_448.fifo_rd_block = 0;
    assign fifo_intf_448.fifo_wr_block = 0;
    assign fifo_intf_448.finish = finish;
    csv_file_dump fifo_csv_dumper_448;
    csv_file_dump cstatus_csv_dumper_448;
    df_fifo_monitor fifo_monitor_448;
    df_fifo_intf fifo_intf_449(clock,reset);
    assign fifo_intf_449.rd_en = AESL_inst_myproject.layer2_out_448_U.if_read & AESL_inst_myproject.layer2_out_448_U.if_empty_n;
    assign fifo_intf_449.wr_en = AESL_inst_myproject.layer2_out_448_U.if_write & AESL_inst_myproject.layer2_out_448_U.if_full_n;
    assign fifo_intf_449.fifo_rd_block = 0;
    assign fifo_intf_449.fifo_wr_block = 0;
    assign fifo_intf_449.finish = finish;
    csv_file_dump fifo_csv_dumper_449;
    csv_file_dump cstatus_csv_dumper_449;
    df_fifo_monitor fifo_monitor_449;
    df_fifo_intf fifo_intf_450(clock,reset);
    assign fifo_intf_450.rd_en = AESL_inst_myproject.layer2_out_449_U.if_read & AESL_inst_myproject.layer2_out_449_U.if_empty_n;
    assign fifo_intf_450.wr_en = AESL_inst_myproject.layer2_out_449_U.if_write & AESL_inst_myproject.layer2_out_449_U.if_full_n;
    assign fifo_intf_450.fifo_rd_block = 0;
    assign fifo_intf_450.fifo_wr_block = 0;
    assign fifo_intf_450.finish = finish;
    csv_file_dump fifo_csv_dumper_450;
    csv_file_dump cstatus_csv_dumper_450;
    df_fifo_monitor fifo_monitor_450;
    df_fifo_intf fifo_intf_451(clock,reset);
    assign fifo_intf_451.rd_en = AESL_inst_myproject.layer2_out_450_U.if_read & AESL_inst_myproject.layer2_out_450_U.if_empty_n;
    assign fifo_intf_451.wr_en = AESL_inst_myproject.layer2_out_450_U.if_write & AESL_inst_myproject.layer2_out_450_U.if_full_n;
    assign fifo_intf_451.fifo_rd_block = 0;
    assign fifo_intf_451.fifo_wr_block = 0;
    assign fifo_intf_451.finish = finish;
    csv_file_dump fifo_csv_dumper_451;
    csv_file_dump cstatus_csv_dumper_451;
    df_fifo_monitor fifo_monitor_451;
    df_fifo_intf fifo_intf_452(clock,reset);
    assign fifo_intf_452.rd_en = AESL_inst_myproject.layer2_out_451_U.if_read & AESL_inst_myproject.layer2_out_451_U.if_empty_n;
    assign fifo_intf_452.wr_en = AESL_inst_myproject.layer2_out_451_U.if_write & AESL_inst_myproject.layer2_out_451_U.if_full_n;
    assign fifo_intf_452.fifo_rd_block = 0;
    assign fifo_intf_452.fifo_wr_block = 0;
    assign fifo_intf_452.finish = finish;
    csv_file_dump fifo_csv_dumper_452;
    csv_file_dump cstatus_csv_dumper_452;
    df_fifo_monitor fifo_monitor_452;
    df_fifo_intf fifo_intf_453(clock,reset);
    assign fifo_intf_453.rd_en = AESL_inst_myproject.layer2_out_452_U.if_read & AESL_inst_myproject.layer2_out_452_U.if_empty_n;
    assign fifo_intf_453.wr_en = AESL_inst_myproject.layer2_out_452_U.if_write & AESL_inst_myproject.layer2_out_452_U.if_full_n;
    assign fifo_intf_453.fifo_rd_block = 0;
    assign fifo_intf_453.fifo_wr_block = 0;
    assign fifo_intf_453.finish = finish;
    csv_file_dump fifo_csv_dumper_453;
    csv_file_dump cstatus_csv_dumper_453;
    df_fifo_monitor fifo_monitor_453;
    df_fifo_intf fifo_intf_454(clock,reset);
    assign fifo_intf_454.rd_en = AESL_inst_myproject.layer2_out_453_U.if_read & AESL_inst_myproject.layer2_out_453_U.if_empty_n;
    assign fifo_intf_454.wr_en = AESL_inst_myproject.layer2_out_453_U.if_write & AESL_inst_myproject.layer2_out_453_U.if_full_n;
    assign fifo_intf_454.fifo_rd_block = 0;
    assign fifo_intf_454.fifo_wr_block = 0;
    assign fifo_intf_454.finish = finish;
    csv_file_dump fifo_csv_dumper_454;
    csv_file_dump cstatus_csv_dumper_454;
    df_fifo_monitor fifo_monitor_454;
    df_fifo_intf fifo_intf_455(clock,reset);
    assign fifo_intf_455.rd_en = AESL_inst_myproject.layer2_out_454_U.if_read & AESL_inst_myproject.layer2_out_454_U.if_empty_n;
    assign fifo_intf_455.wr_en = AESL_inst_myproject.layer2_out_454_U.if_write & AESL_inst_myproject.layer2_out_454_U.if_full_n;
    assign fifo_intf_455.fifo_rd_block = 0;
    assign fifo_intf_455.fifo_wr_block = 0;
    assign fifo_intf_455.finish = finish;
    csv_file_dump fifo_csv_dumper_455;
    csv_file_dump cstatus_csv_dumper_455;
    df_fifo_monitor fifo_monitor_455;
    df_fifo_intf fifo_intf_456(clock,reset);
    assign fifo_intf_456.rd_en = AESL_inst_myproject.layer2_out_455_U.if_read & AESL_inst_myproject.layer2_out_455_U.if_empty_n;
    assign fifo_intf_456.wr_en = AESL_inst_myproject.layer2_out_455_U.if_write & AESL_inst_myproject.layer2_out_455_U.if_full_n;
    assign fifo_intf_456.fifo_rd_block = 0;
    assign fifo_intf_456.fifo_wr_block = 0;
    assign fifo_intf_456.finish = finish;
    csv_file_dump fifo_csv_dumper_456;
    csv_file_dump cstatus_csv_dumper_456;
    df_fifo_monitor fifo_monitor_456;
    df_fifo_intf fifo_intf_457(clock,reset);
    assign fifo_intf_457.rd_en = AESL_inst_myproject.layer2_out_456_U.if_read & AESL_inst_myproject.layer2_out_456_U.if_empty_n;
    assign fifo_intf_457.wr_en = AESL_inst_myproject.layer2_out_456_U.if_write & AESL_inst_myproject.layer2_out_456_U.if_full_n;
    assign fifo_intf_457.fifo_rd_block = 0;
    assign fifo_intf_457.fifo_wr_block = 0;
    assign fifo_intf_457.finish = finish;
    csv_file_dump fifo_csv_dumper_457;
    csv_file_dump cstatus_csv_dumper_457;
    df_fifo_monitor fifo_monitor_457;
    df_fifo_intf fifo_intf_458(clock,reset);
    assign fifo_intf_458.rd_en = AESL_inst_myproject.layer2_out_457_U.if_read & AESL_inst_myproject.layer2_out_457_U.if_empty_n;
    assign fifo_intf_458.wr_en = AESL_inst_myproject.layer2_out_457_U.if_write & AESL_inst_myproject.layer2_out_457_U.if_full_n;
    assign fifo_intf_458.fifo_rd_block = 0;
    assign fifo_intf_458.fifo_wr_block = 0;
    assign fifo_intf_458.finish = finish;
    csv_file_dump fifo_csv_dumper_458;
    csv_file_dump cstatus_csv_dumper_458;
    df_fifo_monitor fifo_monitor_458;
    df_fifo_intf fifo_intf_459(clock,reset);
    assign fifo_intf_459.rd_en = AESL_inst_myproject.layer2_out_458_U.if_read & AESL_inst_myproject.layer2_out_458_U.if_empty_n;
    assign fifo_intf_459.wr_en = AESL_inst_myproject.layer2_out_458_U.if_write & AESL_inst_myproject.layer2_out_458_U.if_full_n;
    assign fifo_intf_459.fifo_rd_block = 0;
    assign fifo_intf_459.fifo_wr_block = 0;
    assign fifo_intf_459.finish = finish;
    csv_file_dump fifo_csv_dumper_459;
    csv_file_dump cstatus_csv_dumper_459;
    df_fifo_monitor fifo_monitor_459;
    df_fifo_intf fifo_intf_460(clock,reset);
    assign fifo_intf_460.rd_en = AESL_inst_myproject.layer2_out_459_U.if_read & AESL_inst_myproject.layer2_out_459_U.if_empty_n;
    assign fifo_intf_460.wr_en = AESL_inst_myproject.layer2_out_459_U.if_write & AESL_inst_myproject.layer2_out_459_U.if_full_n;
    assign fifo_intf_460.fifo_rd_block = 0;
    assign fifo_intf_460.fifo_wr_block = 0;
    assign fifo_intf_460.finish = finish;
    csv_file_dump fifo_csv_dumper_460;
    csv_file_dump cstatus_csv_dumper_460;
    df_fifo_monitor fifo_monitor_460;
    df_fifo_intf fifo_intf_461(clock,reset);
    assign fifo_intf_461.rd_en = AESL_inst_myproject.layer2_out_460_U.if_read & AESL_inst_myproject.layer2_out_460_U.if_empty_n;
    assign fifo_intf_461.wr_en = AESL_inst_myproject.layer2_out_460_U.if_write & AESL_inst_myproject.layer2_out_460_U.if_full_n;
    assign fifo_intf_461.fifo_rd_block = 0;
    assign fifo_intf_461.fifo_wr_block = 0;
    assign fifo_intf_461.finish = finish;
    csv_file_dump fifo_csv_dumper_461;
    csv_file_dump cstatus_csv_dumper_461;
    df_fifo_monitor fifo_monitor_461;
    df_fifo_intf fifo_intf_462(clock,reset);
    assign fifo_intf_462.rd_en = AESL_inst_myproject.layer2_out_461_U.if_read & AESL_inst_myproject.layer2_out_461_U.if_empty_n;
    assign fifo_intf_462.wr_en = AESL_inst_myproject.layer2_out_461_U.if_write & AESL_inst_myproject.layer2_out_461_U.if_full_n;
    assign fifo_intf_462.fifo_rd_block = 0;
    assign fifo_intf_462.fifo_wr_block = 0;
    assign fifo_intf_462.finish = finish;
    csv_file_dump fifo_csv_dumper_462;
    csv_file_dump cstatus_csv_dumper_462;
    df_fifo_monitor fifo_monitor_462;
    df_fifo_intf fifo_intf_463(clock,reset);
    assign fifo_intf_463.rd_en = AESL_inst_myproject.layer2_out_462_U.if_read & AESL_inst_myproject.layer2_out_462_U.if_empty_n;
    assign fifo_intf_463.wr_en = AESL_inst_myproject.layer2_out_462_U.if_write & AESL_inst_myproject.layer2_out_462_U.if_full_n;
    assign fifo_intf_463.fifo_rd_block = 0;
    assign fifo_intf_463.fifo_wr_block = 0;
    assign fifo_intf_463.finish = finish;
    csv_file_dump fifo_csv_dumper_463;
    csv_file_dump cstatus_csv_dumper_463;
    df_fifo_monitor fifo_monitor_463;
    df_fifo_intf fifo_intf_464(clock,reset);
    assign fifo_intf_464.rd_en = AESL_inst_myproject.layer2_out_463_U.if_read & AESL_inst_myproject.layer2_out_463_U.if_empty_n;
    assign fifo_intf_464.wr_en = AESL_inst_myproject.layer2_out_463_U.if_write & AESL_inst_myproject.layer2_out_463_U.if_full_n;
    assign fifo_intf_464.fifo_rd_block = 0;
    assign fifo_intf_464.fifo_wr_block = 0;
    assign fifo_intf_464.finish = finish;
    csv_file_dump fifo_csv_dumper_464;
    csv_file_dump cstatus_csv_dumper_464;
    df_fifo_monitor fifo_monitor_464;
    df_fifo_intf fifo_intf_465(clock,reset);
    assign fifo_intf_465.rd_en = AESL_inst_myproject.layer2_out_464_U.if_read & AESL_inst_myproject.layer2_out_464_U.if_empty_n;
    assign fifo_intf_465.wr_en = AESL_inst_myproject.layer2_out_464_U.if_write & AESL_inst_myproject.layer2_out_464_U.if_full_n;
    assign fifo_intf_465.fifo_rd_block = 0;
    assign fifo_intf_465.fifo_wr_block = 0;
    assign fifo_intf_465.finish = finish;
    csv_file_dump fifo_csv_dumper_465;
    csv_file_dump cstatus_csv_dumper_465;
    df_fifo_monitor fifo_monitor_465;
    df_fifo_intf fifo_intf_466(clock,reset);
    assign fifo_intf_466.rd_en = AESL_inst_myproject.layer2_out_465_U.if_read & AESL_inst_myproject.layer2_out_465_U.if_empty_n;
    assign fifo_intf_466.wr_en = AESL_inst_myproject.layer2_out_465_U.if_write & AESL_inst_myproject.layer2_out_465_U.if_full_n;
    assign fifo_intf_466.fifo_rd_block = 0;
    assign fifo_intf_466.fifo_wr_block = 0;
    assign fifo_intf_466.finish = finish;
    csv_file_dump fifo_csv_dumper_466;
    csv_file_dump cstatus_csv_dumper_466;
    df_fifo_monitor fifo_monitor_466;
    df_fifo_intf fifo_intf_467(clock,reset);
    assign fifo_intf_467.rd_en = AESL_inst_myproject.layer2_out_466_U.if_read & AESL_inst_myproject.layer2_out_466_U.if_empty_n;
    assign fifo_intf_467.wr_en = AESL_inst_myproject.layer2_out_466_U.if_write & AESL_inst_myproject.layer2_out_466_U.if_full_n;
    assign fifo_intf_467.fifo_rd_block = 0;
    assign fifo_intf_467.fifo_wr_block = 0;
    assign fifo_intf_467.finish = finish;
    csv_file_dump fifo_csv_dumper_467;
    csv_file_dump cstatus_csv_dumper_467;
    df_fifo_monitor fifo_monitor_467;
    df_fifo_intf fifo_intf_468(clock,reset);
    assign fifo_intf_468.rd_en = AESL_inst_myproject.layer2_out_467_U.if_read & AESL_inst_myproject.layer2_out_467_U.if_empty_n;
    assign fifo_intf_468.wr_en = AESL_inst_myproject.layer2_out_467_U.if_write & AESL_inst_myproject.layer2_out_467_U.if_full_n;
    assign fifo_intf_468.fifo_rd_block = 0;
    assign fifo_intf_468.fifo_wr_block = 0;
    assign fifo_intf_468.finish = finish;
    csv_file_dump fifo_csv_dumper_468;
    csv_file_dump cstatus_csv_dumper_468;
    df_fifo_monitor fifo_monitor_468;
    df_fifo_intf fifo_intf_469(clock,reset);
    assign fifo_intf_469.rd_en = AESL_inst_myproject.layer2_out_468_U.if_read & AESL_inst_myproject.layer2_out_468_U.if_empty_n;
    assign fifo_intf_469.wr_en = AESL_inst_myproject.layer2_out_468_U.if_write & AESL_inst_myproject.layer2_out_468_U.if_full_n;
    assign fifo_intf_469.fifo_rd_block = 0;
    assign fifo_intf_469.fifo_wr_block = 0;
    assign fifo_intf_469.finish = finish;
    csv_file_dump fifo_csv_dumper_469;
    csv_file_dump cstatus_csv_dumper_469;
    df_fifo_monitor fifo_monitor_469;
    df_fifo_intf fifo_intf_470(clock,reset);
    assign fifo_intf_470.rd_en = AESL_inst_myproject.layer2_out_469_U.if_read & AESL_inst_myproject.layer2_out_469_U.if_empty_n;
    assign fifo_intf_470.wr_en = AESL_inst_myproject.layer2_out_469_U.if_write & AESL_inst_myproject.layer2_out_469_U.if_full_n;
    assign fifo_intf_470.fifo_rd_block = 0;
    assign fifo_intf_470.fifo_wr_block = 0;
    assign fifo_intf_470.finish = finish;
    csv_file_dump fifo_csv_dumper_470;
    csv_file_dump cstatus_csv_dumper_470;
    df_fifo_monitor fifo_monitor_470;
    df_fifo_intf fifo_intf_471(clock,reset);
    assign fifo_intf_471.rd_en = AESL_inst_myproject.layer2_out_470_U.if_read & AESL_inst_myproject.layer2_out_470_U.if_empty_n;
    assign fifo_intf_471.wr_en = AESL_inst_myproject.layer2_out_470_U.if_write & AESL_inst_myproject.layer2_out_470_U.if_full_n;
    assign fifo_intf_471.fifo_rd_block = 0;
    assign fifo_intf_471.fifo_wr_block = 0;
    assign fifo_intf_471.finish = finish;
    csv_file_dump fifo_csv_dumper_471;
    csv_file_dump cstatus_csv_dumper_471;
    df_fifo_monitor fifo_monitor_471;
    df_fifo_intf fifo_intf_472(clock,reset);
    assign fifo_intf_472.rd_en = AESL_inst_myproject.layer2_out_471_U.if_read & AESL_inst_myproject.layer2_out_471_U.if_empty_n;
    assign fifo_intf_472.wr_en = AESL_inst_myproject.layer2_out_471_U.if_write & AESL_inst_myproject.layer2_out_471_U.if_full_n;
    assign fifo_intf_472.fifo_rd_block = 0;
    assign fifo_intf_472.fifo_wr_block = 0;
    assign fifo_intf_472.finish = finish;
    csv_file_dump fifo_csv_dumper_472;
    csv_file_dump cstatus_csv_dumper_472;
    df_fifo_monitor fifo_monitor_472;
    df_fifo_intf fifo_intf_473(clock,reset);
    assign fifo_intf_473.rd_en = AESL_inst_myproject.layer2_out_472_U.if_read & AESL_inst_myproject.layer2_out_472_U.if_empty_n;
    assign fifo_intf_473.wr_en = AESL_inst_myproject.layer2_out_472_U.if_write & AESL_inst_myproject.layer2_out_472_U.if_full_n;
    assign fifo_intf_473.fifo_rd_block = 0;
    assign fifo_intf_473.fifo_wr_block = 0;
    assign fifo_intf_473.finish = finish;
    csv_file_dump fifo_csv_dumper_473;
    csv_file_dump cstatus_csv_dumper_473;
    df_fifo_monitor fifo_monitor_473;
    df_fifo_intf fifo_intf_474(clock,reset);
    assign fifo_intf_474.rd_en = AESL_inst_myproject.layer2_out_473_U.if_read & AESL_inst_myproject.layer2_out_473_U.if_empty_n;
    assign fifo_intf_474.wr_en = AESL_inst_myproject.layer2_out_473_U.if_write & AESL_inst_myproject.layer2_out_473_U.if_full_n;
    assign fifo_intf_474.fifo_rd_block = 0;
    assign fifo_intf_474.fifo_wr_block = 0;
    assign fifo_intf_474.finish = finish;
    csv_file_dump fifo_csv_dumper_474;
    csv_file_dump cstatus_csv_dumper_474;
    df_fifo_monitor fifo_monitor_474;
    df_fifo_intf fifo_intf_475(clock,reset);
    assign fifo_intf_475.rd_en = AESL_inst_myproject.layer2_out_474_U.if_read & AESL_inst_myproject.layer2_out_474_U.if_empty_n;
    assign fifo_intf_475.wr_en = AESL_inst_myproject.layer2_out_474_U.if_write & AESL_inst_myproject.layer2_out_474_U.if_full_n;
    assign fifo_intf_475.fifo_rd_block = 0;
    assign fifo_intf_475.fifo_wr_block = 0;
    assign fifo_intf_475.finish = finish;
    csv_file_dump fifo_csv_dumper_475;
    csv_file_dump cstatus_csv_dumper_475;
    df_fifo_monitor fifo_monitor_475;
    df_fifo_intf fifo_intf_476(clock,reset);
    assign fifo_intf_476.rd_en = AESL_inst_myproject.layer2_out_475_U.if_read & AESL_inst_myproject.layer2_out_475_U.if_empty_n;
    assign fifo_intf_476.wr_en = AESL_inst_myproject.layer2_out_475_U.if_write & AESL_inst_myproject.layer2_out_475_U.if_full_n;
    assign fifo_intf_476.fifo_rd_block = 0;
    assign fifo_intf_476.fifo_wr_block = 0;
    assign fifo_intf_476.finish = finish;
    csv_file_dump fifo_csv_dumper_476;
    csv_file_dump cstatus_csv_dumper_476;
    df_fifo_monitor fifo_monitor_476;
    df_fifo_intf fifo_intf_477(clock,reset);
    assign fifo_intf_477.rd_en = AESL_inst_myproject.layer2_out_476_U.if_read & AESL_inst_myproject.layer2_out_476_U.if_empty_n;
    assign fifo_intf_477.wr_en = AESL_inst_myproject.layer2_out_476_U.if_write & AESL_inst_myproject.layer2_out_476_U.if_full_n;
    assign fifo_intf_477.fifo_rd_block = 0;
    assign fifo_intf_477.fifo_wr_block = 0;
    assign fifo_intf_477.finish = finish;
    csv_file_dump fifo_csv_dumper_477;
    csv_file_dump cstatus_csv_dumper_477;
    df_fifo_monitor fifo_monitor_477;
    df_fifo_intf fifo_intf_478(clock,reset);
    assign fifo_intf_478.rd_en = AESL_inst_myproject.layer2_out_477_U.if_read & AESL_inst_myproject.layer2_out_477_U.if_empty_n;
    assign fifo_intf_478.wr_en = AESL_inst_myproject.layer2_out_477_U.if_write & AESL_inst_myproject.layer2_out_477_U.if_full_n;
    assign fifo_intf_478.fifo_rd_block = 0;
    assign fifo_intf_478.fifo_wr_block = 0;
    assign fifo_intf_478.finish = finish;
    csv_file_dump fifo_csv_dumper_478;
    csv_file_dump cstatus_csv_dumper_478;
    df_fifo_monitor fifo_monitor_478;
    df_fifo_intf fifo_intf_479(clock,reset);
    assign fifo_intf_479.rd_en = AESL_inst_myproject.layer2_out_478_U.if_read & AESL_inst_myproject.layer2_out_478_U.if_empty_n;
    assign fifo_intf_479.wr_en = AESL_inst_myproject.layer2_out_478_U.if_write & AESL_inst_myproject.layer2_out_478_U.if_full_n;
    assign fifo_intf_479.fifo_rd_block = 0;
    assign fifo_intf_479.fifo_wr_block = 0;
    assign fifo_intf_479.finish = finish;
    csv_file_dump fifo_csv_dumper_479;
    csv_file_dump cstatus_csv_dumper_479;
    df_fifo_monitor fifo_monitor_479;
    df_fifo_intf fifo_intf_480(clock,reset);
    assign fifo_intf_480.rd_en = AESL_inst_myproject.layer2_out_479_U.if_read & AESL_inst_myproject.layer2_out_479_U.if_empty_n;
    assign fifo_intf_480.wr_en = AESL_inst_myproject.layer2_out_479_U.if_write & AESL_inst_myproject.layer2_out_479_U.if_full_n;
    assign fifo_intf_480.fifo_rd_block = 0;
    assign fifo_intf_480.fifo_wr_block = 0;
    assign fifo_intf_480.finish = finish;
    csv_file_dump fifo_csv_dumper_480;
    csv_file_dump cstatus_csv_dumper_480;
    df_fifo_monitor fifo_monitor_480;
    df_fifo_intf fifo_intf_481(clock,reset);
    assign fifo_intf_481.rd_en = AESL_inst_myproject.layer2_out_480_U.if_read & AESL_inst_myproject.layer2_out_480_U.if_empty_n;
    assign fifo_intf_481.wr_en = AESL_inst_myproject.layer2_out_480_U.if_write & AESL_inst_myproject.layer2_out_480_U.if_full_n;
    assign fifo_intf_481.fifo_rd_block = 0;
    assign fifo_intf_481.fifo_wr_block = 0;
    assign fifo_intf_481.finish = finish;
    csv_file_dump fifo_csv_dumper_481;
    csv_file_dump cstatus_csv_dumper_481;
    df_fifo_monitor fifo_monitor_481;
    df_fifo_intf fifo_intf_482(clock,reset);
    assign fifo_intf_482.rd_en = AESL_inst_myproject.layer2_out_481_U.if_read & AESL_inst_myproject.layer2_out_481_U.if_empty_n;
    assign fifo_intf_482.wr_en = AESL_inst_myproject.layer2_out_481_U.if_write & AESL_inst_myproject.layer2_out_481_U.if_full_n;
    assign fifo_intf_482.fifo_rd_block = 0;
    assign fifo_intf_482.fifo_wr_block = 0;
    assign fifo_intf_482.finish = finish;
    csv_file_dump fifo_csv_dumper_482;
    csv_file_dump cstatus_csv_dumper_482;
    df_fifo_monitor fifo_monitor_482;
    df_fifo_intf fifo_intf_483(clock,reset);
    assign fifo_intf_483.rd_en = AESL_inst_myproject.layer2_out_482_U.if_read & AESL_inst_myproject.layer2_out_482_U.if_empty_n;
    assign fifo_intf_483.wr_en = AESL_inst_myproject.layer2_out_482_U.if_write & AESL_inst_myproject.layer2_out_482_U.if_full_n;
    assign fifo_intf_483.fifo_rd_block = 0;
    assign fifo_intf_483.fifo_wr_block = 0;
    assign fifo_intf_483.finish = finish;
    csv_file_dump fifo_csv_dumper_483;
    csv_file_dump cstatus_csv_dumper_483;
    df_fifo_monitor fifo_monitor_483;
    df_fifo_intf fifo_intf_484(clock,reset);
    assign fifo_intf_484.rd_en = AESL_inst_myproject.layer2_out_483_U.if_read & AESL_inst_myproject.layer2_out_483_U.if_empty_n;
    assign fifo_intf_484.wr_en = AESL_inst_myproject.layer2_out_483_U.if_write & AESL_inst_myproject.layer2_out_483_U.if_full_n;
    assign fifo_intf_484.fifo_rd_block = 0;
    assign fifo_intf_484.fifo_wr_block = 0;
    assign fifo_intf_484.finish = finish;
    csv_file_dump fifo_csv_dumper_484;
    csv_file_dump cstatus_csv_dumper_484;
    df_fifo_monitor fifo_monitor_484;
    df_fifo_intf fifo_intf_485(clock,reset);
    assign fifo_intf_485.rd_en = AESL_inst_myproject.layer2_out_484_U.if_read & AESL_inst_myproject.layer2_out_484_U.if_empty_n;
    assign fifo_intf_485.wr_en = AESL_inst_myproject.layer2_out_484_U.if_write & AESL_inst_myproject.layer2_out_484_U.if_full_n;
    assign fifo_intf_485.fifo_rd_block = 0;
    assign fifo_intf_485.fifo_wr_block = 0;
    assign fifo_intf_485.finish = finish;
    csv_file_dump fifo_csv_dumper_485;
    csv_file_dump cstatus_csv_dumper_485;
    df_fifo_monitor fifo_monitor_485;
    df_fifo_intf fifo_intf_486(clock,reset);
    assign fifo_intf_486.rd_en = AESL_inst_myproject.layer2_out_485_U.if_read & AESL_inst_myproject.layer2_out_485_U.if_empty_n;
    assign fifo_intf_486.wr_en = AESL_inst_myproject.layer2_out_485_U.if_write & AESL_inst_myproject.layer2_out_485_U.if_full_n;
    assign fifo_intf_486.fifo_rd_block = 0;
    assign fifo_intf_486.fifo_wr_block = 0;
    assign fifo_intf_486.finish = finish;
    csv_file_dump fifo_csv_dumper_486;
    csv_file_dump cstatus_csv_dumper_486;
    df_fifo_monitor fifo_monitor_486;
    df_fifo_intf fifo_intf_487(clock,reset);
    assign fifo_intf_487.rd_en = AESL_inst_myproject.layer2_out_486_U.if_read & AESL_inst_myproject.layer2_out_486_U.if_empty_n;
    assign fifo_intf_487.wr_en = AESL_inst_myproject.layer2_out_486_U.if_write & AESL_inst_myproject.layer2_out_486_U.if_full_n;
    assign fifo_intf_487.fifo_rd_block = 0;
    assign fifo_intf_487.fifo_wr_block = 0;
    assign fifo_intf_487.finish = finish;
    csv_file_dump fifo_csv_dumper_487;
    csv_file_dump cstatus_csv_dumper_487;
    df_fifo_monitor fifo_monitor_487;
    df_fifo_intf fifo_intf_488(clock,reset);
    assign fifo_intf_488.rd_en = AESL_inst_myproject.layer2_out_487_U.if_read & AESL_inst_myproject.layer2_out_487_U.if_empty_n;
    assign fifo_intf_488.wr_en = AESL_inst_myproject.layer2_out_487_U.if_write & AESL_inst_myproject.layer2_out_487_U.if_full_n;
    assign fifo_intf_488.fifo_rd_block = 0;
    assign fifo_intf_488.fifo_wr_block = 0;
    assign fifo_intf_488.finish = finish;
    csv_file_dump fifo_csv_dumper_488;
    csv_file_dump cstatus_csv_dumper_488;
    df_fifo_monitor fifo_monitor_488;
    df_fifo_intf fifo_intf_489(clock,reset);
    assign fifo_intf_489.rd_en = AESL_inst_myproject.layer2_out_488_U.if_read & AESL_inst_myproject.layer2_out_488_U.if_empty_n;
    assign fifo_intf_489.wr_en = AESL_inst_myproject.layer2_out_488_U.if_write & AESL_inst_myproject.layer2_out_488_U.if_full_n;
    assign fifo_intf_489.fifo_rd_block = 0;
    assign fifo_intf_489.fifo_wr_block = 0;
    assign fifo_intf_489.finish = finish;
    csv_file_dump fifo_csv_dumper_489;
    csv_file_dump cstatus_csv_dumper_489;
    df_fifo_monitor fifo_monitor_489;
    df_fifo_intf fifo_intf_490(clock,reset);
    assign fifo_intf_490.rd_en = AESL_inst_myproject.layer2_out_489_U.if_read & AESL_inst_myproject.layer2_out_489_U.if_empty_n;
    assign fifo_intf_490.wr_en = AESL_inst_myproject.layer2_out_489_U.if_write & AESL_inst_myproject.layer2_out_489_U.if_full_n;
    assign fifo_intf_490.fifo_rd_block = 0;
    assign fifo_intf_490.fifo_wr_block = 0;
    assign fifo_intf_490.finish = finish;
    csv_file_dump fifo_csv_dumper_490;
    csv_file_dump cstatus_csv_dumper_490;
    df_fifo_monitor fifo_monitor_490;
    df_fifo_intf fifo_intf_491(clock,reset);
    assign fifo_intf_491.rd_en = AESL_inst_myproject.layer2_out_490_U.if_read & AESL_inst_myproject.layer2_out_490_U.if_empty_n;
    assign fifo_intf_491.wr_en = AESL_inst_myproject.layer2_out_490_U.if_write & AESL_inst_myproject.layer2_out_490_U.if_full_n;
    assign fifo_intf_491.fifo_rd_block = 0;
    assign fifo_intf_491.fifo_wr_block = 0;
    assign fifo_intf_491.finish = finish;
    csv_file_dump fifo_csv_dumper_491;
    csv_file_dump cstatus_csv_dumper_491;
    df_fifo_monitor fifo_monitor_491;
    df_fifo_intf fifo_intf_492(clock,reset);
    assign fifo_intf_492.rd_en = AESL_inst_myproject.layer2_out_491_U.if_read & AESL_inst_myproject.layer2_out_491_U.if_empty_n;
    assign fifo_intf_492.wr_en = AESL_inst_myproject.layer2_out_491_U.if_write & AESL_inst_myproject.layer2_out_491_U.if_full_n;
    assign fifo_intf_492.fifo_rd_block = 0;
    assign fifo_intf_492.fifo_wr_block = 0;
    assign fifo_intf_492.finish = finish;
    csv_file_dump fifo_csv_dumper_492;
    csv_file_dump cstatus_csv_dumper_492;
    df_fifo_monitor fifo_monitor_492;
    df_fifo_intf fifo_intf_493(clock,reset);
    assign fifo_intf_493.rd_en = AESL_inst_myproject.layer2_out_492_U.if_read & AESL_inst_myproject.layer2_out_492_U.if_empty_n;
    assign fifo_intf_493.wr_en = AESL_inst_myproject.layer2_out_492_U.if_write & AESL_inst_myproject.layer2_out_492_U.if_full_n;
    assign fifo_intf_493.fifo_rd_block = 0;
    assign fifo_intf_493.fifo_wr_block = 0;
    assign fifo_intf_493.finish = finish;
    csv_file_dump fifo_csv_dumper_493;
    csv_file_dump cstatus_csv_dumper_493;
    df_fifo_monitor fifo_monitor_493;
    df_fifo_intf fifo_intf_494(clock,reset);
    assign fifo_intf_494.rd_en = AESL_inst_myproject.layer2_out_493_U.if_read & AESL_inst_myproject.layer2_out_493_U.if_empty_n;
    assign fifo_intf_494.wr_en = AESL_inst_myproject.layer2_out_493_U.if_write & AESL_inst_myproject.layer2_out_493_U.if_full_n;
    assign fifo_intf_494.fifo_rd_block = 0;
    assign fifo_intf_494.fifo_wr_block = 0;
    assign fifo_intf_494.finish = finish;
    csv_file_dump fifo_csv_dumper_494;
    csv_file_dump cstatus_csv_dumper_494;
    df_fifo_monitor fifo_monitor_494;
    df_fifo_intf fifo_intf_495(clock,reset);
    assign fifo_intf_495.rd_en = AESL_inst_myproject.layer2_out_494_U.if_read & AESL_inst_myproject.layer2_out_494_U.if_empty_n;
    assign fifo_intf_495.wr_en = AESL_inst_myproject.layer2_out_494_U.if_write & AESL_inst_myproject.layer2_out_494_U.if_full_n;
    assign fifo_intf_495.fifo_rd_block = 0;
    assign fifo_intf_495.fifo_wr_block = 0;
    assign fifo_intf_495.finish = finish;
    csv_file_dump fifo_csv_dumper_495;
    csv_file_dump cstatus_csv_dumper_495;
    df_fifo_monitor fifo_monitor_495;
    df_fifo_intf fifo_intf_496(clock,reset);
    assign fifo_intf_496.rd_en = AESL_inst_myproject.layer2_out_495_U.if_read & AESL_inst_myproject.layer2_out_495_U.if_empty_n;
    assign fifo_intf_496.wr_en = AESL_inst_myproject.layer2_out_495_U.if_write & AESL_inst_myproject.layer2_out_495_U.if_full_n;
    assign fifo_intf_496.fifo_rd_block = 0;
    assign fifo_intf_496.fifo_wr_block = 0;
    assign fifo_intf_496.finish = finish;
    csv_file_dump fifo_csv_dumper_496;
    csv_file_dump cstatus_csv_dumper_496;
    df_fifo_monitor fifo_monitor_496;
    df_fifo_intf fifo_intf_497(clock,reset);
    assign fifo_intf_497.rd_en = AESL_inst_myproject.layer2_out_496_U.if_read & AESL_inst_myproject.layer2_out_496_U.if_empty_n;
    assign fifo_intf_497.wr_en = AESL_inst_myproject.layer2_out_496_U.if_write & AESL_inst_myproject.layer2_out_496_U.if_full_n;
    assign fifo_intf_497.fifo_rd_block = 0;
    assign fifo_intf_497.fifo_wr_block = 0;
    assign fifo_intf_497.finish = finish;
    csv_file_dump fifo_csv_dumper_497;
    csv_file_dump cstatus_csv_dumper_497;
    df_fifo_monitor fifo_monitor_497;
    df_fifo_intf fifo_intf_498(clock,reset);
    assign fifo_intf_498.rd_en = AESL_inst_myproject.layer2_out_497_U.if_read & AESL_inst_myproject.layer2_out_497_U.if_empty_n;
    assign fifo_intf_498.wr_en = AESL_inst_myproject.layer2_out_497_U.if_write & AESL_inst_myproject.layer2_out_497_U.if_full_n;
    assign fifo_intf_498.fifo_rd_block = 0;
    assign fifo_intf_498.fifo_wr_block = 0;
    assign fifo_intf_498.finish = finish;
    csv_file_dump fifo_csv_dumper_498;
    csv_file_dump cstatus_csv_dumper_498;
    df_fifo_monitor fifo_monitor_498;
    df_fifo_intf fifo_intf_499(clock,reset);
    assign fifo_intf_499.rd_en = AESL_inst_myproject.layer2_out_498_U.if_read & AESL_inst_myproject.layer2_out_498_U.if_empty_n;
    assign fifo_intf_499.wr_en = AESL_inst_myproject.layer2_out_498_U.if_write & AESL_inst_myproject.layer2_out_498_U.if_full_n;
    assign fifo_intf_499.fifo_rd_block = 0;
    assign fifo_intf_499.fifo_wr_block = 0;
    assign fifo_intf_499.finish = finish;
    csv_file_dump fifo_csv_dumper_499;
    csv_file_dump cstatus_csv_dumper_499;
    df_fifo_monitor fifo_monitor_499;
    df_fifo_intf fifo_intf_500(clock,reset);
    assign fifo_intf_500.rd_en = AESL_inst_myproject.layer2_out_499_U.if_read & AESL_inst_myproject.layer2_out_499_U.if_empty_n;
    assign fifo_intf_500.wr_en = AESL_inst_myproject.layer2_out_499_U.if_write & AESL_inst_myproject.layer2_out_499_U.if_full_n;
    assign fifo_intf_500.fifo_rd_block = 0;
    assign fifo_intf_500.fifo_wr_block = 0;
    assign fifo_intf_500.finish = finish;
    csv_file_dump fifo_csv_dumper_500;
    csv_file_dump cstatus_csv_dumper_500;
    df_fifo_monitor fifo_monitor_500;
    df_fifo_intf fifo_intf_501(clock,reset);
    assign fifo_intf_501.rd_en = AESL_inst_myproject.layer2_out_500_U.if_read & AESL_inst_myproject.layer2_out_500_U.if_empty_n;
    assign fifo_intf_501.wr_en = AESL_inst_myproject.layer2_out_500_U.if_write & AESL_inst_myproject.layer2_out_500_U.if_full_n;
    assign fifo_intf_501.fifo_rd_block = 0;
    assign fifo_intf_501.fifo_wr_block = 0;
    assign fifo_intf_501.finish = finish;
    csv_file_dump fifo_csv_dumper_501;
    csv_file_dump cstatus_csv_dumper_501;
    df_fifo_monitor fifo_monitor_501;
    df_fifo_intf fifo_intf_502(clock,reset);
    assign fifo_intf_502.rd_en = AESL_inst_myproject.layer2_out_501_U.if_read & AESL_inst_myproject.layer2_out_501_U.if_empty_n;
    assign fifo_intf_502.wr_en = AESL_inst_myproject.layer2_out_501_U.if_write & AESL_inst_myproject.layer2_out_501_U.if_full_n;
    assign fifo_intf_502.fifo_rd_block = 0;
    assign fifo_intf_502.fifo_wr_block = 0;
    assign fifo_intf_502.finish = finish;
    csv_file_dump fifo_csv_dumper_502;
    csv_file_dump cstatus_csv_dumper_502;
    df_fifo_monitor fifo_monitor_502;
    df_fifo_intf fifo_intf_503(clock,reset);
    assign fifo_intf_503.rd_en = AESL_inst_myproject.layer2_out_502_U.if_read & AESL_inst_myproject.layer2_out_502_U.if_empty_n;
    assign fifo_intf_503.wr_en = AESL_inst_myproject.layer2_out_502_U.if_write & AESL_inst_myproject.layer2_out_502_U.if_full_n;
    assign fifo_intf_503.fifo_rd_block = 0;
    assign fifo_intf_503.fifo_wr_block = 0;
    assign fifo_intf_503.finish = finish;
    csv_file_dump fifo_csv_dumper_503;
    csv_file_dump cstatus_csv_dumper_503;
    df_fifo_monitor fifo_monitor_503;
    df_fifo_intf fifo_intf_504(clock,reset);
    assign fifo_intf_504.rd_en = AESL_inst_myproject.layer2_out_503_U.if_read & AESL_inst_myproject.layer2_out_503_U.if_empty_n;
    assign fifo_intf_504.wr_en = AESL_inst_myproject.layer2_out_503_U.if_write & AESL_inst_myproject.layer2_out_503_U.if_full_n;
    assign fifo_intf_504.fifo_rd_block = 0;
    assign fifo_intf_504.fifo_wr_block = 0;
    assign fifo_intf_504.finish = finish;
    csv_file_dump fifo_csv_dumper_504;
    csv_file_dump cstatus_csv_dumper_504;
    df_fifo_monitor fifo_monitor_504;
    df_fifo_intf fifo_intf_505(clock,reset);
    assign fifo_intf_505.rd_en = AESL_inst_myproject.layer2_out_504_U.if_read & AESL_inst_myproject.layer2_out_504_U.if_empty_n;
    assign fifo_intf_505.wr_en = AESL_inst_myproject.layer2_out_504_U.if_write & AESL_inst_myproject.layer2_out_504_U.if_full_n;
    assign fifo_intf_505.fifo_rd_block = 0;
    assign fifo_intf_505.fifo_wr_block = 0;
    assign fifo_intf_505.finish = finish;
    csv_file_dump fifo_csv_dumper_505;
    csv_file_dump cstatus_csv_dumper_505;
    df_fifo_monitor fifo_monitor_505;
    df_fifo_intf fifo_intf_506(clock,reset);
    assign fifo_intf_506.rd_en = AESL_inst_myproject.layer2_out_505_U.if_read & AESL_inst_myproject.layer2_out_505_U.if_empty_n;
    assign fifo_intf_506.wr_en = AESL_inst_myproject.layer2_out_505_U.if_write & AESL_inst_myproject.layer2_out_505_U.if_full_n;
    assign fifo_intf_506.fifo_rd_block = 0;
    assign fifo_intf_506.fifo_wr_block = 0;
    assign fifo_intf_506.finish = finish;
    csv_file_dump fifo_csv_dumper_506;
    csv_file_dump cstatus_csv_dumper_506;
    df_fifo_monitor fifo_monitor_506;
    df_fifo_intf fifo_intf_507(clock,reset);
    assign fifo_intf_507.rd_en = AESL_inst_myproject.layer2_out_506_U.if_read & AESL_inst_myproject.layer2_out_506_U.if_empty_n;
    assign fifo_intf_507.wr_en = AESL_inst_myproject.layer2_out_506_U.if_write & AESL_inst_myproject.layer2_out_506_U.if_full_n;
    assign fifo_intf_507.fifo_rd_block = 0;
    assign fifo_intf_507.fifo_wr_block = 0;
    assign fifo_intf_507.finish = finish;
    csv_file_dump fifo_csv_dumper_507;
    csv_file_dump cstatus_csv_dumper_507;
    df_fifo_monitor fifo_monitor_507;
    df_fifo_intf fifo_intf_508(clock,reset);
    assign fifo_intf_508.rd_en = AESL_inst_myproject.layer2_out_507_U.if_read & AESL_inst_myproject.layer2_out_507_U.if_empty_n;
    assign fifo_intf_508.wr_en = AESL_inst_myproject.layer2_out_507_U.if_write & AESL_inst_myproject.layer2_out_507_U.if_full_n;
    assign fifo_intf_508.fifo_rd_block = 0;
    assign fifo_intf_508.fifo_wr_block = 0;
    assign fifo_intf_508.finish = finish;
    csv_file_dump fifo_csv_dumper_508;
    csv_file_dump cstatus_csv_dumper_508;
    df_fifo_monitor fifo_monitor_508;
    df_fifo_intf fifo_intf_509(clock,reset);
    assign fifo_intf_509.rd_en = AESL_inst_myproject.layer2_out_508_U.if_read & AESL_inst_myproject.layer2_out_508_U.if_empty_n;
    assign fifo_intf_509.wr_en = AESL_inst_myproject.layer2_out_508_U.if_write & AESL_inst_myproject.layer2_out_508_U.if_full_n;
    assign fifo_intf_509.fifo_rd_block = 0;
    assign fifo_intf_509.fifo_wr_block = 0;
    assign fifo_intf_509.finish = finish;
    csv_file_dump fifo_csv_dumper_509;
    csv_file_dump cstatus_csv_dumper_509;
    df_fifo_monitor fifo_monitor_509;
    df_fifo_intf fifo_intf_510(clock,reset);
    assign fifo_intf_510.rd_en = AESL_inst_myproject.layer2_out_509_U.if_read & AESL_inst_myproject.layer2_out_509_U.if_empty_n;
    assign fifo_intf_510.wr_en = AESL_inst_myproject.layer2_out_509_U.if_write & AESL_inst_myproject.layer2_out_509_U.if_full_n;
    assign fifo_intf_510.fifo_rd_block = 0;
    assign fifo_intf_510.fifo_wr_block = 0;
    assign fifo_intf_510.finish = finish;
    csv_file_dump fifo_csv_dumper_510;
    csv_file_dump cstatus_csv_dumper_510;
    df_fifo_monitor fifo_monitor_510;
    df_fifo_intf fifo_intf_511(clock,reset);
    assign fifo_intf_511.rd_en = AESL_inst_myproject.layer2_out_510_U.if_read & AESL_inst_myproject.layer2_out_510_U.if_empty_n;
    assign fifo_intf_511.wr_en = AESL_inst_myproject.layer2_out_510_U.if_write & AESL_inst_myproject.layer2_out_510_U.if_full_n;
    assign fifo_intf_511.fifo_rd_block = 0;
    assign fifo_intf_511.fifo_wr_block = 0;
    assign fifo_intf_511.finish = finish;
    csv_file_dump fifo_csv_dumper_511;
    csv_file_dump cstatus_csv_dumper_511;
    df_fifo_monitor fifo_monitor_511;
    df_fifo_intf fifo_intf_512(clock,reset);
    assign fifo_intf_512.rd_en = AESL_inst_myproject.layer2_out_511_U.if_read & AESL_inst_myproject.layer2_out_511_U.if_empty_n;
    assign fifo_intf_512.wr_en = AESL_inst_myproject.layer2_out_511_U.if_write & AESL_inst_myproject.layer2_out_511_U.if_full_n;
    assign fifo_intf_512.fifo_rd_block = 0;
    assign fifo_intf_512.fifo_wr_block = 0;
    assign fifo_intf_512.finish = finish;
    csv_file_dump fifo_csv_dumper_512;
    csv_file_dump cstatus_csv_dumper_512;
    df_fifo_monitor fifo_monitor_512;
    df_fifo_intf fifo_intf_513(clock,reset);
    assign fifo_intf_513.rd_en = AESL_inst_myproject.layer2_out_512_U.if_read & AESL_inst_myproject.layer2_out_512_U.if_empty_n;
    assign fifo_intf_513.wr_en = AESL_inst_myproject.layer2_out_512_U.if_write & AESL_inst_myproject.layer2_out_512_U.if_full_n;
    assign fifo_intf_513.fifo_rd_block = 0;
    assign fifo_intf_513.fifo_wr_block = 0;
    assign fifo_intf_513.finish = finish;
    csv_file_dump fifo_csv_dumper_513;
    csv_file_dump cstatus_csv_dumper_513;
    df_fifo_monitor fifo_monitor_513;
    df_fifo_intf fifo_intf_514(clock,reset);
    assign fifo_intf_514.rd_en = AESL_inst_myproject.layer2_out_513_U.if_read & AESL_inst_myproject.layer2_out_513_U.if_empty_n;
    assign fifo_intf_514.wr_en = AESL_inst_myproject.layer2_out_513_U.if_write & AESL_inst_myproject.layer2_out_513_U.if_full_n;
    assign fifo_intf_514.fifo_rd_block = 0;
    assign fifo_intf_514.fifo_wr_block = 0;
    assign fifo_intf_514.finish = finish;
    csv_file_dump fifo_csv_dumper_514;
    csv_file_dump cstatus_csv_dumper_514;
    df_fifo_monitor fifo_monitor_514;
    df_fifo_intf fifo_intf_515(clock,reset);
    assign fifo_intf_515.rd_en = AESL_inst_myproject.layer2_out_514_U.if_read & AESL_inst_myproject.layer2_out_514_U.if_empty_n;
    assign fifo_intf_515.wr_en = AESL_inst_myproject.layer2_out_514_U.if_write & AESL_inst_myproject.layer2_out_514_U.if_full_n;
    assign fifo_intf_515.fifo_rd_block = 0;
    assign fifo_intf_515.fifo_wr_block = 0;
    assign fifo_intf_515.finish = finish;
    csv_file_dump fifo_csv_dumper_515;
    csv_file_dump cstatus_csv_dumper_515;
    df_fifo_monitor fifo_monitor_515;
    df_fifo_intf fifo_intf_516(clock,reset);
    assign fifo_intf_516.rd_en = AESL_inst_myproject.layer2_out_515_U.if_read & AESL_inst_myproject.layer2_out_515_U.if_empty_n;
    assign fifo_intf_516.wr_en = AESL_inst_myproject.layer2_out_515_U.if_write & AESL_inst_myproject.layer2_out_515_U.if_full_n;
    assign fifo_intf_516.fifo_rd_block = 0;
    assign fifo_intf_516.fifo_wr_block = 0;
    assign fifo_intf_516.finish = finish;
    csv_file_dump fifo_csv_dumper_516;
    csv_file_dump cstatus_csv_dumper_516;
    df_fifo_monitor fifo_monitor_516;
    df_fifo_intf fifo_intf_517(clock,reset);
    assign fifo_intf_517.rd_en = AESL_inst_myproject.layer2_out_516_U.if_read & AESL_inst_myproject.layer2_out_516_U.if_empty_n;
    assign fifo_intf_517.wr_en = AESL_inst_myproject.layer2_out_516_U.if_write & AESL_inst_myproject.layer2_out_516_U.if_full_n;
    assign fifo_intf_517.fifo_rd_block = 0;
    assign fifo_intf_517.fifo_wr_block = 0;
    assign fifo_intf_517.finish = finish;
    csv_file_dump fifo_csv_dumper_517;
    csv_file_dump cstatus_csv_dumper_517;
    df_fifo_monitor fifo_monitor_517;
    df_fifo_intf fifo_intf_518(clock,reset);
    assign fifo_intf_518.rd_en = AESL_inst_myproject.layer2_out_517_U.if_read & AESL_inst_myproject.layer2_out_517_U.if_empty_n;
    assign fifo_intf_518.wr_en = AESL_inst_myproject.layer2_out_517_U.if_write & AESL_inst_myproject.layer2_out_517_U.if_full_n;
    assign fifo_intf_518.fifo_rd_block = 0;
    assign fifo_intf_518.fifo_wr_block = 0;
    assign fifo_intf_518.finish = finish;
    csv_file_dump fifo_csv_dumper_518;
    csv_file_dump cstatus_csv_dumper_518;
    df_fifo_monitor fifo_monitor_518;
    df_fifo_intf fifo_intf_519(clock,reset);
    assign fifo_intf_519.rd_en = AESL_inst_myproject.layer2_out_518_U.if_read & AESL_inst_myproject.layer2_out_518_U.if_empty_n;
    assign fifo_intf_519.wr_en = AESL_inst_myproject.layer2_out_518_U.if_write & AESL_inst_myproject.layer2_out_518_U.if_full_n;
    assign fifo_intf_519.fifo_rd_block = 0;
    assign fifo_intf_519.fifo_wr_block = 0;
    assign fifo_intf_519.finish = finish;
    csv_file_dump fifo_csv_dumper_519;
    csv_file_dump cstatus_csv_dumper_519;
    df_fifo_monitor fifo_monitor_519;
    df_fifo_intf fifo_intf_520(clock,reset);
    assign fifo_intf_520.rd_en = AESL_inst_myproject.layer2_out_519_U.if_read & AESL_inst_myproject.layer2_out_519_U.if_empty_n;
    assign fifo_intf_520.wr_en = AESL_inst_myproject.layer2_out_519_U.if_write & AESL_inst_myproject.layer2_out_519_U.if_full_n;
    assign fifo_intf_520.fifo_rd_block = 0;
    assign fifo_intf_520.fifo_wr_block = 0;
    assign fifo_intf_520.finish = finish;
    csv_file_dump fifo_csv_dumper_520;
    csv_file_dump cstatus_csv_dumper_520;
    df_fifo_monitor fifo_monitor_520;
    df_fifo_intf fifo_intf_521(clock,reset);
    assign fifo_intf_521.rd_en = AESL_inst_myproject.layer2_out_520_U.if_read & AESL_inst_myproject.layer2_out_520_U.if_empty_n;
    assign fifo_intf_521.wr_en = AESL_inst_myproject.layer2_out_520_U.if_write & AESL_inst_myproject.layer2_out_520_U.if_full_n;
    assign fifo_intf_521.fifo_rd_block = 0;
    assign fifo_intf_521.fifo_wr_block = 0;
    assign fifo_intf_521.finish = finish;
    csv_file_dump fifo_csv_dumper_521;
    csv_file_dump cstatus_csv_dumper_521;
    df_fifo_monitor fifo_monitor_521;
    df_fifo_intf fifo_intf_522(clock,reset);
    assign fifo_intf_522.rd_en = AESL_inst_myproject.layer2_out_521_U.if_read & AESL_inst_myproject.layer2_out_521_U.if_empty_n;
    assign fifo_intf_522.wr_en = AESL_inst_myproject.layer2_out_521_U.if_write & AESL_inst_myproject.layer2_out_521_U.if_full_n;
    assign fifo_intf_522.fifo_rd_block = 0;
    assign fifo_intf_522.fifo_wr_block = 0;
    assign fifo_intf_522.finish = finish;
    csv_file_dump fifo_csv_dumper_522;
    csv_file_dump cstatus_csv_dumper_522;
    df_fifo_monitor fifo_monitor_522;
    df_fifo_intf fifo_intf_523(clock,reset);
    assign fifo_intf_523.rd_en = AESL_inst_myproject.layer2_out_522_U.if_read & AESL_inst_myproject.layer2_out_522_U.if_empty_n;
    assign fifo_intf_523.wr_en = AESL_inst_myproject.layer2_out_522_U.if_write & AESL_inst_myproject.layer2_out_522_U.if_full_n;
    assign fifo_intf_523.fifo_rd_block = 0;
    assign fifo_intf_523.fifo_wr_block = 0;
    assign fifo_intf_523.finish = finish;
    csv_file_dump fifo_csv_dumper_523;
    csv_file_dump cstatus_csv_dumper_523;
    df_fifo_monitor fifo_monitor_523;
    df_fifo_intf fifo_intf_524(clock,reset);
    assign fifo_intf_524.rd_en = AESL_inst_myproject.layer2_out_523_U.if_read & AESL_inst_myproject.layer2_out_523_U.if_empty_n;
    assign fifo_intf_524.wr_en = AESL_inst_myproject.layer2_out_523_U.if_write & AESL_inst_myproject.layer2_out_523_U.if_full_n;
    assign fifo_intf_524.fifo_rd_block = 0;
    assign fifo_intf_524.fifo_wr_block = 0;
    assign fifo_intf_524.finish = finish;
    csv_file_dump fifo_csv_dumper_524;
    csv_file_dump cstatus_csv_dumper_524;
    df_fifo_monitor fifo_monitor_524;
    df_fifo_intf fifo_intf_525(clock,reset);
    assign fifo_intf_525.rd_en = AESL_inst_myproject.layer2_out_524_U.if_read & AESL_inst_myproject.layer2_out_524_U.if_empty_n;
    assign fifo_intf_525.wr_en = AESL_inst_myproject.layer2_out_524_U.if_write & AESL_inst_myproject.layer2_out_524_U.if_full_n;
    assign fifo_intf_525.fifo_rd_block = 0;
    assign fifo_intf_525.fifo_wr_block = 0;
    assign fifo_intf_525.finish = finish;
    csv_file_dump fifo_csv_dumper_525;
    csv_file_dump cstatus_csv_dumper_525;
    df_fifo_monitor fifo_monitor_525;
    df_fifo_intf fifo_intf_526(clock,reset);
    assign fifo_intf_526.rd_en = AESL_inst_myproject.layer2_out_525_U.if_read & AESL_inst_myproject.layer2_out_525_U.if_empty_n;
    assign fifo_intf_526.wr_en = AESL_inst_myproject.layer2_out_525_U.if_write & AESL_inst_myproject.layer2_out_525_U.if_full_n;
    assign fifo_intf_526.fifo_rd_block = 0;
    assign fifo_intf_526.fifo_wr_block = 0;
    assign fifo_intf_526.finish = finish;
    csv_file_dump fifo_csv_dumper_526;
    csv_file_dump cstatus_csv_dumper_526;
    df_fifo_monitor fifo_monitor_526;
    df_fifo_intf fifo_intf_527(clock,reset);
    assign fifo_intf_527.rd_en = AESL_inst_myproject.layer2_out_526_U.if_read & AESL_inst_myproject.layer2_out_526_U.if_empty_n;
    assign fifo_intf_527.wr_en = AESL_inst_myproject.layer2_out_526_U.if_write & AESL_inst_myproject.layer2_out_526_U.if_full_n;
    assign fifo_intf_527.fifo_rd_block = 0;
    assign fifo_intf_527.fifo_wr_block = 0;
    assign fifo_intf_527.finish = finish;
    csv_file_dump fifo_csv_dumper_527;
    csv_file_dump cstatus_csv_dumper_527;
    df_fifo_monitor fifo_monitor_527;
    df_fifo_intf fifo_intf_528(clock,reset);
    assign fifo_intf_528.rd_en = AESL_inst_myproject.layer2_out_527_U.if_read & AESL_inst_myproject.layer2_out_527_U.if_empty_n;
    assign fifo_intf_528.wr_en = AESL_inst_myproject.layer2_out_527_U.if_write & AESL_inst_myproject.layer2_out_527_U.if_full_n;
    assign fifo_intf_528.fifo_rd_block = 0;
    assign fifo_intf_528.fifo_wr_block = 0;
    assign fifo_intf_528.finish = finish;
    csv_file_dump fifo_csv_dumper_528;
    csv_file_dump cstatus_csv_dumper_528;
    df_fifo_monitor fifo_monitor_528;
    df_fifo_intf fifo_intf_529(clock,reset);
    assign fifo_intf_529.rd_en = AESL_inst_myproject.layer2_out_528_U.if_read & AESL_inst_myproject.layer2_out_528_U.if_empty_n;
    assign fifo_intf_529.wr_en = AESL_inst_myproject.layer2_out_528_U.if_write & AESL_inst_myproject.layer2_out_528_U.if_full_n;
    assign fifo_intf_529.fifo_rd_block = 0;
    assign fifo_intf_529.fifo_wr_block = 0;
    assign fifo_intf_529.finish = finish;
    csv_file_dump fifo_csv_dumper_529;
    csv_file_dump cstatus_csv_dumper_529;
    df_fifo_monitor fifo_monitor_529;
    df_fifo_intf fifo_intf_530(clock,reset);
    assign fifo_intf_530.rd_en = AESL_inst_myproject.layer2_out_529_U.if_read & AESL_inst_myproject.layer2_out_529_U.if_empty_n;
    assign fifo_intf_530.wr_en = AESL_inst_myproject.layer2_out_529_U.if_write & AESL_inst_myproject.layer2_out_529_U.if_full_n;
    assign fifo_intf_530.fifo_rd_block = 0;
    assign fifo_intf_530.fifo_wr_block = 0;
    assign fifo_intf_530.finish = finish;
    csv_file_dump fifo_csv_dumper_530;
    csv_file_dump cstatus_csv_dumper_530;
    df_fifo_monitor fifo_monitor_530;
    df_fifo_intf fifo_intf_531(clock,reset);
    assign fifo_intf_531.rd_en = AESL_inst_myproject.layer2_out_530_U.if_read & AESL_inst_myproject.layer2_out_530_U.if_empty_n;
    assign fifo_intf_531.wr_en = AESL_inst_myproject.layer2_out_530_U.if_write & AESL_inst_myproject.layer2_out_530_U.if_full_n;
    assign fifo_intf_531.fifo_rd_block = 0;
    assign fifo_intf_531.fifo_wr_block = 0;
    assign fifo_intf_531.finish = finish;
    csv_file_dump fifo_csv_dumper_531;
    csv_file_dump cstatus_csv_dumper_531;
    df_fifo_monitor fifo_monitor_531;
    df_fifo_intf fifo_intf_532(clock,reset);
    assign fifo_intf_532.rd_en = AESL_inst_myproject.layer2_out_531_U.if_read & AESL_inst_myproject.layer2_out_531_U.if_empty_n;
    assign fifo_intf_532.wr_en = AESL_inst_myproject.layer2_out_531_U.if_write & AESL_inst_myproject.layer2_out_531_U.if_full_n;
    assign fifo_intf_532.fifo_rd_block = 0;
    assign fifo_intf_532.fifo_wr_block = 0;
    assign fifo_intf_532.finish = finish;
    csv_file_dump fifo_csv_dumper_532;
    csv_file_dump cstatus_csv_dumper_532;
    df_fifo_monitor fifo_monitor_532;
    df_fifo_intf fifo_intf_533(clock,reset);
    assign fifo_intf_533.rd_en = AESL_inst_myproject.layer2_out_532_U.if_read & AESL_inst_myproject.layer2_out_532_U.if_empty_n;
    assign fifo_intf_533.wr_en = AESL_inst_myproject.layer2_out_532_U.if_write & AESL_inst_myproject.layer2_out_532_U.if_full_n;
    assign fifo_intf_533.fifo_rd_block = 0;
    assign fifo_intf_533.fifo_wr_block = 0;
    assign fifo_intf_533.finish = finish;
    csv_file_dump fifo_csv_dumper_533;
    csv_file_dump cstatus_csv_dumper_533;
    df_fifo_monitor fifo_monitor_533;
    df_fifo_intf fifo_intf_534(clock,reset);
    assign fifo_intf_534.rd_en = AESL_inst_myproject.layer2_out_533_U.if_read & AESL_inst_myproject.layer2_out_533_U.if_empty_n;
    assign fifo_intf_534.wr_en = AESL_inst_myproject.layer2_out_533_U.if_write & AESL_inst_myproject.layer2_out_533_U.if_full_n;
    assign fifo_intf_534.fifo_rd_block = 0;
    assign fifo_intf_534.fifo_wr_block = 0;
    assign fifo_intf_534.finish = finish;
    csv_file_dump fifo_csv_dumper_534;
    csv_file_dump cstatus_csv_dumper_534;
    df_fifo_monitor fifo_monitor_534;
    df_fifo_intf fifo_intf_535(clock,reset);
    assign fifo_intf_535.rd_en = AESL_inst_myproject.layer2_out_534_U.if_read & AESL_inst_myproject.layer2_out_534_U.if_empty_n;
    assign fifo_intf_535.wr_en = AESL_inst_myproject.layer2_out_534_U.if_write & AESL_inst_myproject.layer2_out_534_U.if_full_n;
    assign fifo_intf_535.fifo_rd_block = 0;
    assign fifo_intf_535.fifo_wr_block = 0;
    assign fifo_intf_535.finish = finish;
    csv_file_dump fifo_csv_dumper_535;
    csv_file_dump cstatus_csv_dumper_535;
    df_fifo_monitor fifo_monitor_535;
    df_fifo_intf fifo_intf_536(clock,reset);
    assign fifo_intf_536.rd_en = AESL_inst_myproject.layer2_out_535_U.if_read & AESL_inst_myproject.layer2_out_535_U.if_empty_n;
    assign fifo_intf_536.wr_en = AESL_inst_myproject.layer2_out_535_U.if_write & AESL_inst_myproject.layer2_out_535_U.if_full_n;
    assign fifo_intf_536.fifo_rd_block = 0;
    assign fifo_intf_536.fifo_wr_block = 0;
    assign fifo_intf_536.finish = finish;
    csv_file_dump fifo_csv_dumper_536;
    csv_file_dump cstatus_csv_dumper_536;
    df_fifo_monitor fifo_monitor_536;
    df_fifo_intf fifo_intf_537(clock,reset);
    assign fifo_intf_537.rd_en = AESL_inst_myproject.layer2_out_536_U.if_read & AESL_inst_myproject.layer2_out_536_U.if_empty_n;
    assign fifo_intf_537.wr_en = AESL_inst_myproject.layer2_out_536_U.if_write & AESL_inst_myproject.layer2_out_536_U.if_full_n;
    assign fifo_intf_537.fifo_rd_block = 0;
    assign fifo_intf_537.fifo_wr_block = 0;
    assign fifo_intf_537.finish = finish;
    csv_file_dump fifo_csv_dumper_537;
    csv_file_dump cstatus_csv_dumper_537;
    df_fifo_monitor fifo_monitor_537;
    df_fifo_intf fifo_intf_538(clock,reset);
    assign fifo_intf_538.rd_en = AESL_inst_myproject.layer2_out_537_U.if_read & AESL_inst_myproject.layer2_out_537_U.if_empty_n;
    assign fifo_intf_538.wr_en = AESL_inst_myproject.layer2_out_537_U.if_write & AESL_inst_myproject.layer2_out_537_U.if_full_n;
    assign fifo_intf_538.fifo_rd_block = 0;
    assign fifo_intf_538.fifo_wr_block = 0;
    assign fifo_intf_538.finish = finish;
    csv_file_dump fifo_csv_dumper_538;
    csv_file_dump cstatus_csv_dumper_538;
    df_fifo_monitor fifo_monitor_538;
    df_fifo_intf fifo_intf_539(clock,reset);
    assign fifo_intf_539.rd_en = AESL_inst_myproject.layer2_out_538_U.if_read & AESL_inst_myproject.layer2_out_538_U.if_empty_n;
    assign fifo_intf_539.wr_en = AESL_inst_myproject.layer2_out_538_U.if_write & AESL_inst_myproject.layer2_out_538_U.if_full_n;
    assign fifo_intf_539.fifo_rd_block = 0;
    assign fifo_intf_539.fifo_wr_block = 0;
    assign fifo_intf_539.finish = finish;
    csv_file_dump fifo_csv_dumper_539;
    csv_file_dump cstatus_csv_dumper_539;
    df_fifo_monitor fifo_monitor_539;
    df_fifo_intf fifo_intf_540(clock,reset);
    assign fifo_intf_540.rd_en = AESL_inst_myproject.layer2_out_539_U.if_read & AESL_inst_myproject.layer2_out_539_U.if_empty_n;
    assign fifo_intf_540.wr_en = AESL_inst_myproject.layer2_out_539_U.if_write & AESL_inst_myproject.layer2_out_539_U.if_full_n;
    assign fifo_intf_540.fifo_rd_block = 0;
    assign fifo_intf_540.fifo_wr_block = 0;
    assign fifo_intf_540.finish = finish;
    csv_file_dump fifo_csv_dumper_540;
    csv_file_dump cstatus_csv_dumper_540;
    df_fifo_monitor fifo_monitor_540;
    df_fifo_intf fifo_intf_541(clock,reset);
    assign fifo_intf_541.rd_en = AESL_inst_myproject.layer2_out_540_U.if_read & AESL_inst_myproject.layer2_out_540_U.if_empty_n;
    assign fifo_intf_541.wr_en = AESL_inst_myproject.layer2_out_540_U.if_write & AESL_inst_myproject.layer2_out_540_U.if_full_n;
    assign fifo_intf_541.fifo_rd_block = 0;
    assign fifo_intf_541.fifo_wr_block = 0;
    assign fifo_intf_541.finish = finish;
    csv_file_dump fifo_csv_dumper_541;
    csv_file_dump cstatus_csv_dumper_541;
    df_fifo_monitor fifo_monitor_541;
    df_fifo_intf fifo_intf_542(clock,reset);
    assign fifo_intf_542.rd_en = AESL_inst_myproject.layer2_out_541_U.if_read & AESL_inst_myproject.layer2_out_541_U.if_empty_n;
    assign fifo_intf_542.wr_en = AESL_inst_myproject.layer2_out_541_U.if_write & AESL_inst_myproject.layer2_out_541_U.if_full_n;
    assign fifo_intf_542.fifo_rd_block = 0;
    assign fifo_intf_542.fifo_wr_block = 0;
    assign fifo_intf_542.finish = finish;
    csv_file_dump fifo_csv_dumper_542;
    csv_file_dump cstatus_csv_dumper_542;
    df_fifo_monitor fifo_monitor_542;
    df_fifo_intf fifo_intf_543(clock,reset);
    assign fifo_intf_543.rd_en = AESL_inst_myproject.layer2_out_542_U.if_read & AESL_inst_myproject.layer2_out_542_U.if_empty_n;
    assign fifo_intf_543.wr_en = AESL_inst_myproject.layer2_out_542_U.if_write & AESL_inst_myproject.layer2_out_542_U.if_full_n;
    assign fifo_intf_543.fifo_rd_block = 0;
    assign fifo_intf_543.fifo_wr_block = 0;
    assign fifo_intf_543.finish = finish;
    csv_file_dump fifo_csv_dumper_543;
    csv_file_dump cstatus_csv_dumper_543;
    df_fifo_monitor fifo_monitor_543;
    df_fifo_intf fifo_intf_544(clock,reset);
    assign fifo_intf_544.rd_en = AESL_inst_myproject.layer2_out_543_U.if_read & AESL_inst_myproject.layer2_out_543_U.if_empty_n;
    assign fifo_intf_544.wr_en = AESL_inst_myproject.layer2_out_543_U.if_write & AESL_inst_myproject.layer2_out_543_U.if_full_n;
    assign fifo_intf_544.fifo_rd_block = 0;
    assign fifo_intf_544.fifo_wr_block = 0;
    assign fifo_intf_544.finish = finish;
    csv_file_dump fifo_csv_dumper_544;
    csv_file_dump cstatus_csv_dumper_544;
    df_fifo_monitor fifo_monitor_544;
    df_fifo_intf fifo_intf_545(clock,reset);
    assign fifo_intf_545.rd_en = AESL_inst_myproject.layer2_out_544_U.if_read & AESL_inst_myproject.layer2_out_544_U.if_empty_n;
    assign fifo_intf_545.wr_en = AESL_inst_myproject.layer2_out_544_U.if_write & AESL_inst_myproject.layer2_out_544_U.if_full_n;
    assign fifo_intf_545.fifo_rd_block = 0;
    assign fifo_intf_545.fifo_wr_block = 0;
    assign fifo_intf_545.finish = finish;
    csv_file_dump fifo_csv_dumper_545;
    csv_file_dump cstatus_csv_dumper_545;
    df_fifo_monitor fifo_monitor_545;
    df_fifo_intf fifo_intf_546(clock,reset);
    assign fifo_intf_546.rd_en = AESL_inst_myproject.layer2_out_545_U.if_read & AESL_inst_myproject.layer2_out_545_U.if_empty_n;
    assign fifo_intf_546.wr_en = AESL_inst_myproject.layer2_out_545_U.if_write & AESL_inst_myproject.layer2_out_545_U.if_full_n;
    assign fifo_intf_546.fifo_rd_block = 0;
    assign fifo_intf_546.fifo_wr_block = 0;
    assign fifo_intf_546.finish = finish;
    csv_file_dump fifo_csv_dumper_546;
    csv_file_dump cstatus_csv_dumper_546;
    df_fifo_monitor fifo_monitor_546;
    df_fifo_intf fifo_intf_547(clock,reset);
    assign fifo_intf_547.rd_en = AESL_inst_myproject.layer2_out_546_U.if_read & AESL_inst_myproject.layer2_out_546_U.if_empty_n;
    assign fifo_intf_547.wr_en = AESL_inst_myproject.layer2_out_546_U.if_write & AESL_inst_myproject.layer2_out_546_U.if_full_n;
    assign fifo_intf_547.fifo_rd_block = 0;
    assign fifo_intf_547.fifo_wr_block = 0;
    assign fifo_intf_547.finish = finish;
    csv_file_dump fifo_csv_dumper_547;
    csv_file_dump cstatus_csv_dumper_547;
    df_fifo_monitor fifo_monitor_547;
    df_fifo_intf fifo_intf_548(clock,reset);
    assign fifo_intf_548.rd_en = AESL_inst_myproject.layer2_out_547_U.if_read & AESL_inst_myproject.layer2_out_547_U.if_empty_n;
    assign fifo_intf_548.wr_en = AESL_inst_myproject.layer2_out_547_U.if_write & AESL_inst_myproject.layer2_out_547_U.if_full_n;
    assign fifo_intf_548.fifo_rd_block = 0;
    assign fifo_intf_548.fifo_wr_block = 0;
    assign fifo_intf_548.finish = finish;
    csv_file_dump fifo_csv_dumper_548;
    csv_file_dump cstatus_csv_dumper_548;
    df_fifo_monitor fifo_monitor_548;
    df_fifo_intf fifo_intf_549(clock,reset);
    assign fifo_intf_549.rd_en = AESL_inst_myproject.layer2_out_548_U.if_read & AESL_inst_myproject.layer2_out_548_U.if_empty_n;
    assign fifo_intf_549.wr_en = AESL_inst_myproject.layer2_out_548_U.if_write & AESL_inst_myproject.layer2_out_548_U.if_full_n;
    assign fifo_intf_549.fifo_rd_block = 0;
    assign fifo_intf_549.fifo_wr_block = 0;
    assign fifo_intf_549.finish = finish;
    csv_file_dump fifo_csv_dumper_549;
    csv_file_dump cstatus_csv_dumper_549;
    df_fifo_monitor fifo_monitor_549;
    df_fifo_intf fifo_intf_550(clock,reset);
    assign fifo_intf_550.rd_en = AESL_inst_myproject.layer2_out_549_U.if_read & AESL_inst_myproject.layer2_out_549_U.if_empty_n;
    assign fifo_intf_550.wr_en = AESL_inst_myproject.layer2_out_549_U.if_write & AESL_inst_myproject.layer2_out_549_U.if_full_n;
    assign fifo_intf_550.fifo_rd_block = 0;
    assign fifo_intf_550.fifo_wr_block = 0;
    assign fifo_intf_550.finish = finish;
    csv_file_dump fifo_csv_dumper_550;
    csv_file_dump cstatus_csv_dumper_550;
    df_fifo_monitor fifo_monitor_550;
    df_fifo_intf fifo_intf_551(clock,reset);
    assign fifo_intf_551.rd_en = AESL_inst_myproject.layer2_out_550_U.if_read & AESL_inst_myproject.layer2_out_550_U.if_empty_n;
    assign fifo_intf_551.wr_en = AESL_inst_myproject.layer2_out_550_U.if_write & AESL_inst_myproject.layer2_out_550_U.if_full_n;
    assign fifo_intf_551.fifo_rd_block = 0;
    assign fifo_intf_551.fifo_wr_block = 0;
    assign fifo_intf_551.finish = finish;
    csv_file_dump fifo_csv_dumper_551;
    csv_file_dump cstatus_csv_dumper_551;
    df_fifo_monitor fifo_monitor_551;
    df_fifo_intf fifo_intf_552(clock,reset);
    assign fifo_intf_552.rd_en = AESL_inst_myproject.layer2_out_551_U.if_read & AESL_inst_myproject.layer2_out_551_U.if_empty_n;
    assign fifo_intf_552.wr_en = AESL_inst_myproject.layer2_out_551_U.if_write & AESL_inst_myproject.layer2_out_551_U.if_full_n;
    assign fifo_intf_552.fifo_rd_block = 0;
    assign fifo_intf_552.fifo_wr_block = 0;
    assign fifo_intf_552.finish = finish;
    csv_file_dump fifo_csv_dumper_552;
    csv_file_dump cstatus_csv_dumper_552;
    df_fifo_monitor fifo_monitor_552;
    df_fifo_intf fifo_intf_553(clock,reset);
    assign fifo_intf_553.rd_en = AESL_inst_myproject.layer2_out_552_U.if_read & AESL_inst_myproject.layer2_out_552_U.if_empty_n;
    assign fifo_intf_553.wr_en = AESL_inst_myproject.layer2_out_552_U.if_write & AESL_inst_myproject.layer2_out_552_U.if_full_n;
    assign fifo_intf_553.fifo_rd_block = 0;
    assign fifo_intf_553.fifo_wr_block = 0;
    assign fifo_intf_553.finish = finish;
    csv_file_dump fifo_csv_dumper_553;
    csv_file_dump cstatus_csv_dumper_553;
    df_fifo_monitor fifo_monitor_553;
    df_fifo_intf fifo_intf_554(clock,reset);
    assign fifo_intf_554.rd_en = AESL_inst_myproject.layer2_out_553_U.if_read & AESL_inst_myproject.layer2_out_553_U.if_empty_n;
    assign fifo_intf_554.wr_en = AESL_inst_myproject.layer2_out_553_U.if_write & AESL_inst_myproject.layer2_out_553_U.if_full_n;
    assign fifo_intf_554.fifo_rd_block = 0;
    assign fifo_intf_554.fifo_wr_block = 0;
    assign fifo_intf_554.finish = finish;
    csv_file_dump fifo_csv_dumper_554;
    csv_file_dump cstatus_csv_dumper_554;
    df_fifo_monitor fifo_monitor_554;
    df_fifo_intf fifo_intf_555(clock,reset);
    assign fifo_intf_555.rd_en = AESL_inst_myproject.layer2_out_554_U.if_read & AESL_inst_myproject.layer2_out_554_U.if_empty_n;
    assign fifo_intf_555.wr_en = AESL_inst_myproject.layer2_out_554_U.if_write & AESL_inst_myproject.layer2_out_554_U.if_full_n;
    assign fifo_intf_555.fifo_rd_block = 0;
    assign fifo_intf_555.fifo_wr_block = 0;
    assign fifo_intf_555.finish = finish;
    csv_file_dump fifo_csv_dumper_555;
    csv_file_dump cstatus_csv_dumper_555;
    df_fifo_monitor fifo_monitor_555;
    df_fifo_intf fifo_intf_556(clock,reset);
    assign fifo_intf_556.rd_en = AESL_inst_myproject.layer2_out_555_U.if_read & AESL_inst_myproject.layer2_out_555_U.if_empty_n;
    assign fifo_intf_556.wr_en = AESL_inst_myproject.layer2_out_555_U.if_write & AESL_inst_myproject.layer2_out_555_U.if_full_n;
    assign fifo_intf_556.fifo_rd_block = 0;
    assign fifo_intf_556.fifo_wr_block = 0;
    assign fifo_intf_556.finish = finish;
    csv_file_dump fifo_csv_dumper_556;
    csv_file_dump cstatus_csv_dumper_556;
    df_fifo_monitor fifo_monitor_556;
    df_fifo_intf fifo_intf_557(clock,reset);
    assign fifo_intf_557.rd_en = AESL_inst_myproject.layer2_out_556_U.if_read & AESL_inst_myproject.layer2_out_556_U.if_empty_n;
    assign fifo_intf_557.wr_en = AESL_inst_myproject.layer2_out_556_U.if_write & AESL_inst_myproject.layer2_out_556_U.if_full_n;
    assign fifo_intf_557.fifo_rd_block = 0;
    assign fifo_intf_557.fifo_wr_block = 0;
    assign fifo_intf_557.finish = finish;
    csv_file_dump fifo_csv_dumper_557;
    csv_file_dump cstatus_csv_dumper_557;
    df_fifo_monitor fifo_monitor_557;
    df_fifo_intf fifo_intf_558(clock,reset);
    assign fifo_intf_558.rd_en = AESL_inst_myproject.layer2_out_557_U.if_read & AESL_inst_myproject.layer2_out_557_U.if_empty_n;
    assign fifo_intf_558.wr_en = AESL_inst_myproject.layer2_out_557_U.if_write & AESL_inst_myproject.layer2_out_557_U.if_full_n;
    assign fifo_intf_558.fifo_rd_block = 0;
    assign fifo_intf_558.fifo_wr_block = 0;
    assign fifo_intf_558.finish = finish;
    csv_file_dump fifo_csv_dumper_558;
    csv_file_dump cstatus_csv_dumper_558;
    df_fifo_monitor fifo_monitor_558;
    df_fifo_intf fifo_intf_559(clock,reset);
    assign fifo_intf_559.rd_en = AESL_inst_myproject.layer2_out_558_U.if_read & AESL_inst_myproject.layer2_out_558_U.if_empty_n;
    assign fifo_intf_559.wr_en = AESL_inst_myproject.layer2_out_558_U.if_write & AESL_inst_myproject.layer2_out_558_U.if_full_n;
    assign fifo_intf_559.fifo_rd_block = 0;
    assign fifo_intf_559.fifo_wr_block = 0;
    assign fifo_intf_559.finish = finish;
    csv_file_dump fifo_csv_dumper_559;
    csv_file_dump cstatus_csv_dumper_559;
    df_fifo_monitor fifo_monitor_559;
    df_fifo_intf fifo_intf_560(clock,reset);
    assign fifo_intf_560.rd_en = AESL_inst_myproject.layer2_out_559_U.if_read & AESL_inst_myproject.layer2_out_559_U.if_empty_n;
    assign fifo_intf_560.wr_en = AESL_inst_myproject.layer2_out_559_U.if_write & AESL_inst_myproject.layer2_out_559_U.if_full_n;
    assign fifo_intf_560.fifo_rd_block = 0;
    assign fifo_intf_560.fifo_wr_block = 0;
    assign fifo_intf_560.finish = finish;
    csv_file_dump fifo_csv_dumper_560;
    csv_file_dump cstatus_csv_dumper_560;
    df_fifo_monitor fifo_monitor_560;
    df_fifo_intf fifo_intf_561(clock,reset);
    assign fifo_intf_561.rd_en = AESL_inst_myproject.layer2_out_560_U.if_read & AESL_inst_myproject.layer2_out_560_U.if_empty_n;
    assign fifo_intf_561.wr_en = AESL_inst_myproject.layer2_out_560_U.if_write & AESL_inst_myproject.layer2_out_560_U.if_full_n;
    assign fifo_intf_561.fifo_rd_block = 0;
    assign fifo_intf_561.fifo_wr_block = 0;
    assign fifo_intf_561.finish = finish;
    csv_file_dump fifo_csv_dumper_561;
    csv_file_dump cstatus_csv_dumper_561;
    df_fifo_monitor fifo_monitor_561;
    df_fifo_intf fifo_intf_562(clock,reset);
    assign fifo_intf_562.rd_en = AESL_inst_myproject.layer2_out_561_U.if_read & AESL_inst_myproject.layer2_out_561_U.if_empty_n;
    assign fifo_intf_562.wr_en = AESL_inst_myproject.layer2_out_561_U.if_write & AESL_inst_myproject.layer2_out_561_U.if_full_n;
    assign fifo_intf_562.fifo_rd_block = 0;
    assign fifo_intf_562.fifo_wr_block = 0;
    assign fifo_intf_562.finish = finish;
    csv_file_dump fifo_csv_dumper_562;
    csv_file_dump cstatus_csv_dumper_562;
    df_fifo_monitor fifo_monitor_562;
    df_fifo_intf fifo_intf_563(clock,reset);
    assign fifo_intf_563.rd_en = AESL_inst_myproject.layer2_out_562_U.if_read & AESL_inst_myproject.layer2_out_562_U.if_empty_n;
    assign fifo_intf_563.wr_en = AESL_inst_myproject.layer2_out_562_U.if_write & AESL_inst_myproject.layer2_out_562_U.if_full_n;
    assign fifo_intf_563.fifo_rd_block = 0;
    assign fifo_intf_563.fifo_wr_block = 0;
    assign fifo_intf_563.finish = finish;
    csv_file_dump fifo_csv_dumper_563;
    csv_file_dump cstatus_csv_dumper_563;
    df_fifo_monitor fifo_monitor_563;
    df_fifo_intf fifo_intf_564(clock,reset);
    assign fifo_intf_564.rd_en = AESL_inst_myproject.layer2_out_563_U.if_read & AESL_inst_myproject.layer2_out_563_U.if_empty_n;
    assign fifo_intf_564.wr_en = AESL_inst_myproject.layer2_out_563_U.if_write & AESL_inst_myproject.layer2_out_563_U.if_full_n;
    assign fifo_intf_564.fifo_rd_block = 0;
    assign fifo_intf_564.fifo_wr_block = 0;
    assign fifo_intf_564.finish = finish;
    csv_file_dump fifo_csv_dumper_564;
    csv_file_dump cstatus_csv_dumper_564;
    df_fifo_monitor fifo_monitor_564;
    df_fifo_intf fifo_intf_565(clock,reset);
    assign fifo_intf_565.rd_en = AESL_inst_myproject.layer2_out_564_U.if_read & AESL_inst_myproject.layer2_out_564_U.if_empty_n;
    assign fifo_intf_565.wr_en = AESL_inst_myproject.layer2_out_564_U.if_write & AESL_inst_myproject.layer2_out_564_U.if_full_n;
    assign fifo_intf_565.fifo_rd_block = 0;
    assign fifo_intf_565.fifo_wr_block = 0;
    assign fifo_intf_565.finish = finish;
    csv_file_dump fifo_csv_dumper_565;
    csv_file_dump cstatus_csv_dumper_565;
    df_fifo_monitor fifo_monitor_565;
    df_fifo_intf fifo_intf_566(clock,reset);
    assign fifo_intf_566.rd_en = AESL_inst_myproject.layer2_out_565_U.if_read & AESL_inst_myproject.layer2_out_565_U.if_empty_n;
    assign fifo_intf_566.wr_en = AESL_inst_myproject.layer2_out_565_U.if_write & AESL_inst_myproject.layer2_out_565_U.if_full_n;
    assign fifo_intf_566.fifo_rd_block = 0;
    assign fifo_intf_566.fifo_wr_block = 0;
    assign fifo_intf_566.finish = finish;
    csv_file_dump fifo_csv_dumper_566;
    csv_file_dump cstatus_csv_dumper_566;
    df_fifo_monitor fifo_monitor_566;
    df_fifo_intf fifo_intf_567(clock,reset);
    assign fifo_intf_567.rd_en = AESL_inst_myproject.layer2_out_566_U.if_read & AESL_inst_myproject.layer2_out_566_U.if_empty_n;
    assign fifo_intf_567.wr_en = AESL_inst_myproject.layer2_out_566_U.if_write & AESL_inst_myproject.layer2_out_566_U.if_full_n;
    assign fifo_intf_567.fifo_rd_block = 0;
    assign fifo_intf_567.fifo_wr_block = 0;
    assign fifo_intf_567.finish = finish;
    csv_file_dump fifo_csv_dumper_567;
    csv_file_dump cstatus_csv_dumper_567;
    df_fifo_monitor fifo_monitor_567;
    df_fifo_intf fifo_intf_568(clock,reset);
    assign fifo_intf_568.rd_en = AESL_inst_myproject.layer2_out_567_U.if_read & AESL_inst_myproject.layer2_out_567_U.if_empty_n;
    assign fifo_intf_568.wr_en = AESL_inst_myproject.layer2_out_567_U.if_write & AESL_inst_myproject.layer2_out_567_U.if_full_n;
    assign fifo_intf_568.fifo_rd_block = 0;
    assign fifo_intf_568.fifo_wr_block = 0;
    assign fifo_intf_568.finish = finish;
    csv_file_dump fifo_csv_dumper_568;
    csv_file_dump cstatus_csv_dumper_568;
    df_fifo_monitor fifo_monitor_568;
    df_fifo_intf fifo_intf_569(clock,reset);
    assign fifo_intf_569.rd_en = AESL_inst_myproject.layer2_out_568_U.if_read & AESL_inst_myproject.layer2_out_568_U.if_empty_n;
    assign fifo_intf_569.wr_en = AESL_inst_myproject.layer2_out_568_U.if_write & AESL_inst_myproject.layer2_out_568_U.if_full_n;
    assign fifo_intf_569.fifo_rd_block = 0;
    assign fifo_intf_569.fifo_wr_block = 0;
    assign fifo_intf_569.finish = finish;
    csv_file_dump fifo_csv_dumper_569;
    csv_file_dump cstatus_csv_dumper_569;
    df_fifo_monitor fifo_monitor_569;
    df_fifo_intf fifo_intf_570(clock,reset);
    assign fifo_intf_570.rd_en = AESL_inst_myproject.layer2_out_569_U.if_read & AESL_inst_myproject.layer2_out_569_U.if_empty_n;
    assign fifo_intf_570.wr_en = AESL_inst_myproject.layer2_out_569_U.if_write & AESL_inst_myproject.layer2_out_569_U.if_full_n;
    assign fifo_intf_570.fifo_rd_block = 0;
    assign fifo_intf_570.fifo_wr_block = 0;
    assign fifo_intf_570.finish = finish;
    csv_file_dump fifo_csv_dumper_570;
    csv_file_dump cstatus_csv_dumper_570;
    df_fifo_monitor fifo_monitor_570;
    df_fifo_intf fifo_intf_571(clock,reset);
    assign fifo_intf_571.rd_en = AESL_inst_myproject.layer2_out_570_U.if_read & AESL_inst_myproject.layer2_out_570_U.if_empty_n;
    assign fifo_intf_571.wr_en = AESL_inst_myproject.layer2_out_570_U.if_write & AESL_inst_myproject.layer2_out_570_U.if_full_n;
    assign fifo_intf_571.fifo_rd_block = 0;
    assign fifo_intf_571.fifo_wr_block = 0;
    assign fifo_intf_571.finish = finish;
    csv_file_dump fifo_csv_dumper_571;
    csv_file_dump cstatus_csv_dumper_571;
    df_fifo_monitor fifo_monitor_571;
    df_fifo_intf fifo_intf_572(clock,reset);
    assign fifo_intf_572.rd_en = AESL_inst_myproject.layer2_out_571_U.if_read & AESL_inst_myproject.layer2_out_571_U.if_empty_n;
    assign fifo_intf_572.wr_en = AESL_inst_myproject.layer2_out_571_U.if_write & AESL_inst_myproject.layer2_out_571_U.if_full_n;
    assign fifo_intf_572.fifo_rd_block = 0;
    assign fifo_intf_572.fifo_wr_block = 0;
    assign fifo_intf_572.finish = finish;
    csv_file_dump fifo_csv_dumper_572;
    csv_file_dump cstatus_csv_dumper_572;
    df_fifo_monitor fifo_monitor_572;
    df_fifo_intf fifo_intf_573(clock,reset);
    assign fifo_intf_573.rd_en = AESL_inst_myproject.layer2_out_572_U.if_read & AESL_inst_myproject.layer2_out_572_U.if_empty_n;
    assign fifo_intf_573.wr_en = AESL_inst_myproject.layer2_out_572_U.if_write & AESL_inst_myproject.layer2_out_572_U.if_full_n;
    assign fifo_intf_573.fifo_rd_block = 0;
    assign fifo_intf_573.fifo_wr_block = 0;
    assign fifo_intf_573.finish = finish;
    csv_file_dump fifo_csv_dumper_573;
    csv_file_dump cstatus_csv_dumper_573;
    df_fifo_monitor fifo_monitor_573;
    df_fifo_intf fifo_intf_574(clock,reset);
    assign fifo_intf_574.rd_en = AESL_inst_myproject.layer2_out_573_U.if_read & AESL_inst_myproject.layer2_out_573_U.if_empty_n;
    assign fifo_intf_574.wr_en = AESL_inst_myproject.layer2_out_573_U.if_write & AESL_inst_myproject.layer2_out_573_U.if_full_n;
    assign fifo_intf_574.fifo_rd_block = 0;
    assign fifo_intf_574.fifo_wr_block = 0;
    assign fifo_intf_574.finish = finish;
    csv_file_dump fifo_csv_dumper_574;
    csv_file_dump cstatus_csv_dumper_574;
    df_fifo_monitor fifo_monitor_574;
    df_fifo_intf fifo_intf_575(clock,reset);
    assign fifo_intf_575.rd_en = AESL_inst_myproject.layer2_out_574_U.if_read & AESL_inst_myproject.layer2_out_574_U.if_empty_n;
    assign fifo_intf_575.wr_en = AESL_inst_myproject.layer2_out_574_U.if_write & AESL_inst_myproject.layer2_out_574_U.if_full_n;
    assign fifo_intf_575.fifo_rd_block = 0;
    assign fifo_intf_575.fifo_wr_block = 0;
    assign fifo_intf_575.finish = finish;
    csv_file_dump fifo_csv_dumper_575;
    csv_file_dump cstatus_csv_dumper_575;
    df_fifo_monitor fifo_monitor_575;
    df_fifo_intf fifo_intf_576(clock,reset);
    assign fifo_intf_576.rd_en = AESL_inst_myproject.layer2_out_575_U.if_read & AESL_inst_myproject.layer2_out_575_U.if_empty_n;
    assign fifo_intf_576.wr_en = AESL_inst_myproject.layer2_out_575_U.if_write & AESL_inst_myproject.layer2_out_575_U.if_full_n;
    assign fifo_intf_576.fifo_rd_block = 0;
    assign fifo_intf_576.fifo_wr_block = 0;
    assign fifo_intf_576.finish = finish;
    csv_file_dump fifo_csv_dumper_576;
    csv_file_dump cstatus_csv_dumper_576;
    df_fifo_monitor fifo_monitor_576;
    df_fifo_intf fifo_intf_577(clock,reset);
    assign fifo_intf_577.rd_en = AESL_inst_myproject.layer2_out_576_U.if_read & AESL_inst_myproject.layer2_out_576_U.if_empty_n;
    assign fifo_intf_577.wr_en = AESL_inst_myproject.layer2_out_576_U.if_write & AESL_inst_myproject.layer2_out_576_U.if_full_n;
    assign fifo_intf_577.fifo_rd_block = 0;
    assign fifo_intf_577.fifo_wr_block = 0;
    assign fifo_intf_577.finish = finish;
    csv_file_dump fifo_csv_dumper_577;
    csv_file_dump cstatus_csv_dumper_577;
    df_fifo_monitor fifo_monitor_577;
    df_fifo_intf fifo_intf_578(clock,reset);
    assign fifo_intf_578.rd_en = AESL_inst_myproject.layer2_out_577_U.if_read & AESL_inst_myproject.layer2_out_577_U.if_empty_n;
    assign fifo_intf_578.wr_en = AESL_inst_myproject.layer2_out_577_U.if_write & AESL_inst_myproject.layer2_out_577_U.if_full_n;
    assign fifo_intf_578.fifo_rd_block = 0;
    assign fifo_intf_578.fifo_wr_block = 0;
    assign fifo_intf_578.finish = finish;
    csv_file_dump fifo_csv_dumper_578;
    csv_file_dump cstatus_csv_dumper_578;
    df_fifo_monitor fifo_monitor_578;
    df_fifo_intf fifo_intf_579(clock,reset);
    assign fifo_intf_579.rd_en = AESL_inst_myproject.layer2_out_578_U.if_read & AESL_inst_myproject.layer2_out_578_U.if_empty_n;
    assign fifo_intf_579.wr_en = AESL_inst_myproject.layer2_out_578_U.if_write & AESL_inst_myproject.layer2_out_578_U.if_full_n;
    assign fifo_intf_579.fifo_rd_block = 0;
    assign fifo_intf_579.fifo_wr_block = 0;
    assign fifo_intf_579.finish = finish;
    csv_file_dump fifo_csv_dumper_579;
    csv_file_dump cstatus_csv_dumper_579;
    df_fifo_monitor fifo_monitor_579;
    df_fifo_intf fifo_intf_580(clock,reset);
    assign fifo_intf_580.rd_en = AESL_inst_myproject.layer2_out_579_U.if_read & AESL_inst_myproject.layer2_out_579_U.if_empty_n;
    assign fifo_intf_580.wr_en = AESL_inst_myproject.layer2_out_579_U.if_write & AESL_inst_myproject.layer2_out_579_U.if_full_n;
    assign fifo_intf_580.fifo_rd_block = 0;
    assign fifo_intf_580.fifo_wr_block = 0;
    assign fifo_intf_580.finish = finish;
    csv_file_dump fifo_csv_dumper_580;
    csv_file_dump cstatus_csv_dumper_580;
    df_fifo_monitor fifo_monitor_580;
    df_fifo_intf fifo_intf_581(clock,reset);
    assign fifo_intf_581.rd_en = AESL_inst_myproject.layer2_out_580_U.if_read & AESL_inst_myproject.layer2_out_580_U.if_empty_n;
    assign fifo_intf_581.wr_en = AESL_inst_myproject.layer2_out_580_U.if_write & AESL_inst_myproject.layer2_out_580_U.if_full_n;
    assign fifo_intf_581.fifo_rd_block = 0;
    assign fifo_intf_581.fifo_wr_block = 0;
    assign fifo_intf_581.finish = finish;
    csv_file_dump fifo_csv_dumper_581;
    csv_file_dump cstatus_csv_dumper_581;
    df_fifo_monitor fifo_monitor_581;
    df_fifo_intf fifo_intf_582(clock,reset);
    assign fifo_intf_582.rd_en = AESL_inst_myproject.layer2_out_581_U.if_read & AESL_inst_myproject.layer2_out_581_U.if_empty_n;
    assign fifo_intf_582.wr_en = AESL_inst_myproject.layer2_out_581_U.if_write & AESL_inst_myproject.layer2_out_581_U.if_full_n;
    assign fifo_intf_582.fifo_rd_block = 0;
    assign fifo_intf_582.fifo_wr_block = 0;
    assign fifo_intf_582.finish = finish;
    csv_file_dump fifo_csv_dumper_582;
    csv_file_dump cstatus_csv_dumper_582;
    df_fifo_monitor fifo_monitor_582;
    df_fifo_intf fifo_intf_583(clock,reset);
    assign fifo_intf_583.rd_en = AESL_inst_myproject.layer2_out_582_U.if_read & AESL_inst_myproject.layer2_out_582_U.if_empty_n;
    assign fifo_intf_583.wr_en = AESL_inst_myproject.layer2_out_582_U.if_write & AESL_inst_myproject.layer2_out_582_U.if_full_n;
    assign fifo_intf_583.fifo_rd_block = 0;
    assign fifo_intf_583.fifo_wr_block = 0;
    assign fifo_intf_583.finish = finish;
    csv_file_dump fifo_csv_dumper_583;
    csv_file_dump cstatus_csv_dumper_583;
    df_fifo_monitor fifo_monitor_583;
    df_fifo_intf fifo_intf_584(clock,reset);
    assign fifo_intf_584.rd_en = AESL_inst_myproject.layer2_out_583_U.if_read & AESL_inst_myproject.layer2_out_583_U.if_empty_n;
    assign fifo_intf_584.wr_en = AESL_inst_myproject.layer2_out_583_U.if_write & AESL_inst_myproject.layer2_out_583_U.if_full_n;
    assign fifo_intf_584.fifo_rd_block = 0;
    assign fifo_intf_584.fifo_wr_block = 0;
    assign fifo_intf_584.finish = finish;
    csv_file_dump fifo_csv_dumper_584;
    csv_file_dump cstatus_csv_dumper_584;
    df_fifo_monitor fifo_monitor_584;
    df_fifo_intf fifo_intf_585(clock,reset);
    assign fifo_intf_585.rd_en = AESL_inst_myproject.layer2_out_584_U.if_read & AESL_inst_myproject.layer2_out_584_U.if_empty_n;
    assign fifo_intf_585.wr_en = AESL_inst_myproject.layer2_out_584_U.if_write & AESL_inst_myproject.layer2_out_584_U.if_full_n;
    assign fifo_intf_585.fifo_rd_block = 0;
    assign fifo_intf_585.fifo_wr_block = 0;
    assign fifo_intf_585.finish = finish;
    csv_file_dump fifo_csv_dumper_585;
    csv_file_dump cstatus_csv_dumper_585;
    df_fifo_monitor fifo_monitor_585;
    df_fifo_intf fifo_intf_586(clock,reset);
    assign fifo_intf_586.rd_en = AESL_inst_myproject.layer2_out_585_U.if_read & AESL_inst_myproject.layer2_out_585_U.if_empty_n;
    assign fifo_intf_586.wr_en = AESL_inst_myproject.layer2_out_585_U.if_write & AESL_inst_myproject.layer2_out_585_U.if_full_n;
    assign fifo_intf_586.fifo_rd_block = 0;
    assign fifo_intf_586.fifo_wr_block = 0;
    assign fifo_intf_586.finish = finish;
    csv_file_dump fifo_csv_dumper_586;
    csv_file_dump cstatus_csv_dumper_586;
    df_fifo_monitor fifo_monitor_586;
    df_fifo_intf fifo_intf_587(clock,reset);
    assign fifo_intf_587.rd_en = AESL_inst_myproject.layer2_out_586_U.if_read & AESL_inst_myproject.layer2_out_586_U.if_empty_n;
    assign fifo_intf_587.wr_en = AESL_inst_myproject.layer2_out_586_U.if_write & AESL_inst_myproject.layer2_out_586_U.if_full_n;
    assign fifo_intf_587.fifo_rd_block = 0;
    assign fifo_intf_587.fifo_wr_block = 0;
    assign fifo_intf_587.finish = finish;
    csv_file_dump fifo_csv_dumper_587;
    csv_file_dump cstatus_csv_dumper_587;
    df_fifo_monitor fifo_monitor_587;
    df_fifo_intf fifo_intf_588(clock,reset);
    assign fifo_intf_588.rd_en = AESL_inst_myproject.layer2_out_587_U.if_read & AESL_inst_myproject.layer2_out_587_U.if_empty_n;
    assign fifo_intf_588.wr_en = AESL_inst_myproject.layer2_out_587_U.if_write & AESL_inst_myproject.layer2_out_587_U.if_full_n;
    assign fifo_intf_588.fifo_rd_block = 0;
    assign fifo_intf_588.fifo_wr_block = 0;
    assign fifo_intf_588.finish = finish;
    csv_file_dump fifo_csv_dumper_588;
    csv_file_dump cstatus_csv_dumper_588;
    df_fifo_monitor fifo_monitor_588;
    df_fifo_intf fifo_intf_589(clock,reset);
    assign fifo_intf_589.rd_en = AESL_inst_myproject.layer2_out_588_U.if_read & AESL_inst_myproject.layer2_out_588_U.if_empty_n;
    assign fifo_intf_589.wr_en = AESL_inst_myproject.layer2_out_588_U.if_write & AESL_inst_myproject.layer2_out_588_U.if_full_n;
    assign fifo_intf_589.fifo_rd_block = 0;
    assign fifo_intf_589.fifo_wr_block = 0;
    assign fifo_intf_589.finish = finish;
    csv_file_dump fifo_csv_dumper_589;
    csv_file_dump cstatus_csv_dumper_589;
    df_fifo_monitor fifo_monitor_589;
    df_fifo_intf fifo_intf_590(clock,reset);
    assign fifo_intf_590.rd_en = AESL_inst_myproject.layer2_out_589_U.if_read & AESL_inst_myproject.layer2_out_589_U.if_empty_n;
    assign fifo_intf_590.wr_en = AESL_inst_myproject.layer2_out_589_U.if_write & AESL_inst_myproject.layer2_out_589_U.if_full_n;
    assign fifo_intf_590.fifo_rd_block = 0;
    assign fifo_intf_590.fifo_wr_block = 0;
    assign fifo_intf_590.finish = finish;
    csv_file_dump fifo_csv_dumper_590;
    csv_file_dump cstatus_csv_dumper_590;
    df_fifo_monitor fifo_monitor_590;
    df_fifo_intf fifo_intf_591(clock,reset);
    assign fifo_intf_591.rd_en = AESL_inst_myproject.layer2_out_590_U.if_read & AESL_inst_myproject.layer2_out_590_U.if_empty_n;
    assign fifo_intf_591.wr_en = AESL_inst_myproject.layer2_out_590_U.if_write & AESL_inst_myproject.layer2_out_590_U.if_full_n;
    assign fifo_intf_591.fifo_rd_block = 0;
    assign fifo_intf_591.fifo_wr_block = 0;
    assign fifo_intf_591.finish = finish;
    csv_file_dump fifo_csv_dumper_591;
    csv_file_dump cstatus_csv_dumper_591;
    df_fifo_monitor fifo_monitor_591;
    df_fifo_intf fifo_intf_592(clock,reset);
    assign fifo_intf_592.rd_en = AESL_inst_myproject.layer2_out_591_U.if_read & AESL_inst_myproject.layer2_out_591_U.if_empty_n;
    assign fifo_intf_592.wr_en = AESL_inst_myproject.layer2_out_591_U.if_write & AESL_inst_myproject.layer2_out_591_U.if_full_n;
    assign fifo_intf_592.fifo_rd_block = 0;
    assign fifo_intf_592.fifo_wr_block = 0;
    assign fifo_intf_592.finish = finish;
    csv_file_dump fifo_csv_dumper_592;
    csv_file_dump cstatus_csv_dumper_592;
    df_fifo_monitor fifo_monitor_592;
    df_fifo_intf fifo_intf_593(clock,reset);
    assign fifo_intf_593.rd_en = AESL_inst_myproject.layer2_out_592_U.if_read & AESL_inst_myproject.layer2_out_592_U.if_empty_n;
    assign fifo_intf_593.wr_en = AESL_inst_myproject.layer2_out_592_U.if_write & AESL_inst_myproject.layer2_out_592_U.if_full_n;
    assign fifo_intf_593.fifo_rd_block = 0;
    assign fifo_intf_593.fifo_wr_block = 0;
    assign fifo_intf_593.finish = finish;
    csv_file_dump fifo_csv_dumper_593;
    csv_file_dump cstatus_csv_dumper_593;
    df_fifo_monitor fifo_monitor_593;
    df_fifo_intf fifo_intf_594(clock,reset);
    assign fifo_intf_594.rd_en = AESL_inst_myproject.layer2_out_593_U.if_read & AESL_inst_myproject.layer2_out_593_U.if_empty_n;
    assign fifo_intf_594.wr_en = AESL_inst_myproject.layer2_out_593_U.if_write & AESL_inst_myproject.layer2_out_593_U.if_full_n;
    assign fifo_intf_594.fifo_rd_block = 0;
    assign fifo_intf_594.fifo_wr_block = 0;
    assign fifo_intf_594.finish = finish;
    csv_file_dump fifo_csv_dumper_594;
    csv_file_dump cstatus_csv_dumper_594;
    df_fifo_monitor fifo_monitor_594;
    df_fifo_intf fifo_intf_595(clock,reset);
    assign fifo_intf_595.rd_en = AESL_inst_myproject.layer2_out_594_U.if_read & AESL_inst_myproject.layer2_out_594_U.if_empty_n;
    assign fifo_intf_595.wr_en = AESL_inst_myproject.layer2_out_594_U.if_write & AESL_inst_myproject.layer2_out_594_U.if_full_n;
    assign fifo_intf_595.fifo_rd_block = 0;
    assign fifo_intf_595.fifo_wr_block = 0;
    assign fifo_intf_595.finish = finish;
    csv_file_dump fifo_csv_dumper_595;
    csv_file_dump cstatus_csv_dumper_595;
    df_fifo_monitor fifo_monitor_595;
    df_fifo_intf fifo_intf_596(clock,reset);
    assign fifo_intf_596.rd_en = AESL_inst_myproject.layer2_out_595_U.if_read & AESL_inst_myproject.layer2_out_595_U.if_empty_n;
    assign fifo_intf_596.wr_en = AESL_inst_myproject.layer2_out_595_U.if_write & AESL_inst_myproject.layer2_out_595_U.if_full_n;
    assign fifo_intf_596.fifo_rd_block = 0;
    assign fifo_intf_596.fifo_wr_block = 0;
    assign fifo_intf_596.finish = finish;
    csv_file_dump fifo_csv_dumper_596;
    csv_file_dump cstatus_csv_dumper_596;
    df_fifo_monitor fifo_monitor_596;
    df_fifo_intf fifo_intf_597(clock,reset);
    assign fifo_intf_597.rd_en = AESL_inst_myproject.layer2_out_596_U.if_read & AESL_inst_myproject.layer2_out_596_U.if_empty_n;
    assign fifo_intf_597.wr_en = AESL_inst_myproject.layer2_out_596_U.if_write & AESL_inst_myproject.layer2_out_596_U.if_full_n;
    assign fifo_intf_597.fifo_rd_block = 0;
    assign fifo_intf_597.fifo_wr_block = 0;
    assign fifo_intf_597.finish = finish;
    csv_file_dump fifo_csv_dumper_597;
    csv_file_dump cstatus_csv_dumper_597;
    df_fifo_monitor fifo_monitor_597;
    df_fifo_intf fifo_intf_598(clock,reset);
    assign fifo_intf_598.rd_en = AESL_inst_myproject.layer2_out_597_U.if_read & AESL_inst_myproject.layer2_out_597_U.if_empty_n;
    assign fifo_intf_598.wr_en = AESL_inst_myproject.layer2_out_597_U.if_write & AESL_inst_myproject.layer2_out_597_U.if_full_n;
    assign fifo_intf_598.fifo_rd_block = 0;
    assign fifo_intf_598.fifo_wr_block = 0;
    assign fifo_intf_598.finish = finish;
    csv_file_dump fifo_csv_dumper_598;
    csv_file_dump cstatus_csv_dumper_598;
    df_fifo_monitor fifo_monitor_598;
    df_fifo_intf fifo_intf_599(clock,reset);
    assign fifo_intf_599.rd_en = AESL_inst_myproject.layer2_out_598_U.if_read & AESL_inst_myproject.layer2_out_598_U.if_empty_n;
    assign fifo_intf_599.wr_en = AESL_inst_myproject.layer2_out_598_U.if_write & AESL_inst_myproject.layer2_out_598_U.if_full_n;
    assign fifo_intf_599.fifo_rd_block = 0;
    assign fifo_intf_599.fifo_wr_block = 0;
    assign fifo_intf_599.finish = finish;
    csv_file_dump fifo_csv_dumper_599;
    csv_file_dump cstatus_csv_dumper_599;
    df_fifo_monitor fifo_monitor_599;
    df_fifo_intf fifo_intf_600(clock,reset);
    assign fifo_intf_600.rd_en = AESL_inst_myproject.layer2_out_599_U.if_read & AESL_inst_myproject.layer2_out_599_U.if_empty_n;
    assign fifo_intf_600.wr_en = AESL_inst_myproject.layer2_out_599_U.if_write & AESL_inst_myproject.layer2_out_599_U.if_full_n;
    assign fifo_intf_600.fifo_rd_block = 0;
    assign fifo_intf_600.fifo_wr_block = 0;
    assign fifo_intf_600.finish = finish;
    csv_file_dump fifo_csv_dumper_600;
    csv_file_dump cstatus_csv_dumper_600;
    df_fifo_monitor fifo_monitor_600;
    df_fifo_intf fifo_intf_601(clock,reset);
    assign fifo_intf_601.rd_en = AESL_inst_myproject.layer2_out_600_U.if_read & AESL_inst_myproject.layer2_out_600_U.if_empty_n;
    assign fifo_intf_601.wr_en = AESL_inst_myproject.layer2_out_600_U.if_write & AESL_inst_myproject.layer2_out_600_U.if_full_n;
    assign fifo_intf_601.fifo_rd_block = 0;
    assign fifo_intf_601.fifo_wr_block = 0;
    assign fifo_intf_601.finish = finish;
    csv_file_dump fifo_csv_dumper_601;
    csv_file_dump cstatus_csv_dumper_601;
    df_fifo_monitor fifo_monitor_601;
    df_fifo_intf fifo_intf_602(clock,reset);
    assign fifo_intf_602.rd_en = AESL_inst_myproject.layer2_out_601_U.if_read & AESL_inst_myproject.layer2_out_601_U.if_empty_n;
    assign fifo_intf_602.wr_en = AESL_inst_myproject.layer2_out_601_U.if_write & AESL_inst_myproject.layer2_out_601_U.if_full_n;
    assign fifo_intf_602.fifo_rd_block = 0;
    assign fifo_intf_602.fifo_wr_block = 0;
    assign fifo_intf_602.finish = finish;
    csv_file_dump fifo_csv_dumper_602;
    csv_file_dump cstatus_csv_dumper_602;
    df_fifo_monitor fifo_monitor_602;
    df_fifo_intf fifo_intf_603(clock,reset);
    assign fifo_intf_603.rd_en = AESL_inst_myproject.layer2_out_602_U.if_read & AESL_inst_myproject.layer2_out_602_U.if_empty_n;
    assign fifo_intf_603.wr_en = AESL_inst_myproject.layer2_out_602_U.if_write & AESL_inst_myproject.layer2_out_602_U.if_full_n;
    assign fifo_intf_603.fifo_rd_block = 0;
    assign fifo_intf_603.fifo_wr_block = 0;
    assign fifo_intf_603.finish = finish;
    csv_file_dump fifo_csv_dumper_603;
    csv_file_dump cstatus_csv_dumper_603;
    df_fifo_monitor fifo_monitor_603;
    df_fifo_intf fifo_intf_604(clock,reset);
    assign fifo_intf_604.rd_en = AESL_inst_myproject.layer2_out_603_U.if_read & AESL_inst_myproject.layer2_out_603_U.if_empty_n;
    assign fifo_intf_604.wr_en = AESL_inst_myproject.layer2_out_603_U.if_write & AESL_inst_myproject.layer2_out_603_U.if_full_n;
    assign fifo_intf_604.fifo_rd_block = 0;
    assign fifo_intf_604.fifo_wr_block = 0;
    assign fifo_intf_604.finish = finish;
    csv_file_dump fifo_csv_dumper_604;
    csv_file_dump cstatus_csv_dumper_604;
    df_fifo_monitor fifo_monitor_604;
    df_fifo_intf fifo_intf_605(clock,reset);
    assign fifo_intf_605.rd_en = AESL_inst_myproject.layer2_out_604_U.if_read & AESL_inst_myproject.layer2_out_604_U.if_empty_n;
    assign fifo_intf_605.wr_en = AESL_inst_myproject.layer2_out_604_U.if_write & AESL_inst_myproject.layer2_out_604_U.if_full_n;
    assign fifo_intf_605.fifo_rd_block = 0;
    assign fifo_intf_605.fifo_wr_block = 0;
    assign fifo_intf_605.finish = finish;
    csv_file_dump fifo_csv_dumper_605;
    csv_file_dump cstatus_csv_dumper_605;
    df_fifo_monitor fifo_monitor_605;
    df_fifo_intf fifo_intf_606(clock,reset);
    assign fifo_intf_606.rd_en = AESL_inst_myproject.layer2_out_605_U.if_read & AESL_inst_myproject.layer2_out_605_U.if_empty_n;
    assign fifo_intf_606.wr_en = AESL_inst_myproject.layer2_out_605_U.if_write & AESL_inst_myproject.layer2_out_605_U.if_full_n;
    assign fifo_intf_606.fifo_rd_block = 0;
    assign fifo_intf_606.fifo_wr_block = 0;
    assign fifo_intf_606.finish = finish;
    csv_file_dump fifo_csv_dumper_606;
    csv_file_dump cstatus_csv_dumper_606;
    df_fifo_monitor fifo_monitor_606;
    df_fifo_intf fifo_intf_607(clock,reset);
    assign fifo_intf_607.rd_en = AESL_inst_myproject.layer2_out_606_U.if_read & AESL_inst_myproject.layer2_out_606_U.if_empty_n;
    assign fifo_intf_607.wr_en = AESL_inst_myproject.layer2_out_606_U.if_write & AESL_inst_myproject.layer2_out_606_U.if_full_n;
    assign fifo_intf_607.fifo_rd_block = 0;
    assign fifo_intf_607.fifo_wr_block = 0;
    assign fifo_intf_607.finish = finish;
    csv_file_dump fifo_csv_dumper_607;
    csv_file_dump cstatus_csv_dumper_607;
    df_fifo_monitor fifo_monitor_607;
    df_fifo_intf fifo_intf_608(clock,reset);
    assign fifo_intf_608.rd_en = AESL_inst_myproject.layer2_out_607_U.if_read & AESL_inst_myproject.layer2_out_607_U.if_empty_n;
    assign fifo_intf_608.wr_en = AESL_inst_myproject.layer2_out_607_U.if_write & AESL_inst_myproject.layer2_out_607_U.if_full_n;
    assign fifo_intf_608.fifo_rd_block = 0;
    assign fifo_intf_608.fifo_wr_block = 0;
    assign fifo_intf_608.finish = finish;
    csv_file_dump fifo_csv_dumper_608;
    csv_file_dump cstatus_csv_dumper_608;
    df_fifo_monitor fifo_monitor_608;
    df_fifo_intf fifo_intf_609(clock,reset);
    assign fifo_intf_609.rd_en = AESL_inst_myproject.layer2_out_608_U.if_read & AESL_inst_myproject.layer2_out_608_U.if_empty_n;
    assign fifo_intf_609.wr_en = AESL_inst_myproject.layer2_out_608_U.if_write & AESL_inst_myproject.layer2_out_608_U.if_full_n;
    assign fifo_intf_609.fifo_rd_block = 0;
    assign fifo_intf_609.fifo_wr_block = 0;
    assign fifo_intf_609.finish = finish;
    csv_file_dump fifo_csv_dumper_609;
    csv_file_dump cstatus_csv_dumper_609;
    df_fifo_monitor fifo_monitor_609;
    df_fifo_intf fifo_intf_610(clock,reset);
    assign fifo_intf_610.rd_en = AESL_inst_myproject.layer2_out_609_U.if_read & AESL_inst_myproject.layer2_out_609_U.if_empty_n;
    assign fifo_intf_610.wr_en = AESL_inst_myproject.layer2_out_609_U.if_write & AESL_inst_myproject.layer2_out_609_U.if_full_n;
    assign fifo_intf_610.fifo_rd_block = 0;
    assign fifo_intf_610.fifo_wr_block = 0;
    assign fifo_intf_610.finish = finish;
    csv_file_dump fifo_csv_dumper_610;
    csv_file_dump cstatus_csv_dumper_610;
    df_fifo_monitor fifo_monitor_610;
    df_fifo_intf fifo_intf_611(clock,reset);
    assign fifo_intf_611.rd_en = AESL_inst_myproject.layer2_out_610_U.if_read & AESL_inst_myproject.layer2_out_610_U.if_empty_n;
    assign fifo_intf_611.wr_en = AESL_inst_myproject.layer2_out_610_U.if_write & AESL_inst_myproject.layer2_out_610_U.if_full_n;
    assign fifo_intf_611.fifo_rd_block = 0;
    assign fifo_intf_611.fifo_wr_block = 0;
    assign fifo_intf_611.finish = finish;
    csv_file_dump fifo_csv_dumper_611;
    csv_file_dump cstatus_csv_dumper_611;
    df_fifo_monitor fifo_monitor_611;
    df_fifo_intf fifo_intf_612(clock,reset);
    assign fifo_intf_612.rd_en = AESL_inst_myproject.layer2_out_611_U.if_read & AESL_inst_myproject.layer2_out_611_U.if_empty_n;
    assign fifo_intf_612.wr_en = AESL_inst_myproject.layer2_out_611_U.if_write & AESL_inst_myproject.layer2_out_611_U.if_full_n;
    assign fifo_intf_612.fifo_rd_block = 0;
    assign fifo_intf_612.fifo_wr_block = 0;
    assign fifo_intf_612.finish = finish;
    csv_file_dump fifo_csv_dumper_612;
    csv_file_dump cstatus_csv_dumper_612;
    df_fifo_monitor fifo_monitor_612;
    df_fifo_intf fifo_intf_613(clock,reset);
    assign fifo_intf_613.rd_en = AESL_inst_myproject.layer2_out_612_U.if_read & AESL_inst_myproject.layer2_out_612_U.if_empty_n;
    assign fifo_intf_613.wr_en = AESL_inst_myproject.layer2_out_612_U.if_write & AESL_inst_myproject.layer2_out_612_U.if_full_n;
    assign fifo_intf_613.fifo_rd_block = 0;
    assign fifo_intf_613.fifo_wr_block = 0;
    assign fifo_intf_613.finish = finish;
    csv_file_dump fifo_csv_dumper_613;
    csv_file_dump cstatus_csv_dumper_613;
    df_fifo_monitor fifo_monitor_613;
    df_fifo_intf fifo_intf_614(clock,reset);
    assign fifo_intf_614.rd_en = AESL_inst_myproject.layer2_out_613_U.if_read & AESL_inst_myproject.layer2_out_613_U.if_empty_n;
    assign fifo_intf_614.wr_en = AESL_inst_myproject.layer2_out_613_U.if_write & AESL_inst_myproject.layer2_out_613_U.if_full_n;
    assign fifo_intf_614.fifo_rd_block = 0;
    assign fifo_intf_614.fifo_wr_block = 0;
    assign fifo_intf_614.finish = finish;
    csv_file_dump fifo_csv_dumper_614;
    csv_file_dump cstatus_csv_dumper_614;
    df_fifo_monitor fifo_monitor_614;
    df_fifo_intf fifo_intf_615(clock,reset);
    assign fifo_intf_615.rd_en = AESL_inst_myproject.layer2_out_614_U.if_read & AESL_inst_myproject.layer2_out_614_U.if_empty_n;
    assign fifo_intf_615.wr_en = AESL_inst_myproject.layer2_out_614_U.if_write & AESL_inst_myproject.layer2_out_614_U.if_full_n;
    assign fifo_intf_615.fifo_rd_block = 0;
    assign fifo_intf_615.fifo_wr_block = 0;
    assign fifo_intf_615.finish = finish;
    csv_file_dump fifo_csv_dumper_615;
    csv_file_dump cstatus_csv_dumper_615;
    df_fifo_monitor fifo_monitor_615;
    df_fifo_intf fifo_intf_616(clock,reset);
    assign fifo_intf_616.rd_en = AESL_inst_myproject.layer2_out_615_U.if_read & AESL_inst_myproject.layer2_out_615_U.if_empty_n;
    assign fifo_intf_616.wr_en = AESL_inst_myproject.layer2_out_615_U.if_write & AESL_inst_myproject.layer2_out_615_U.if_full_n;
    assign fifo_intf_616.fifo_rd_block = 0;
    assign fifo_intf_616.fifo_wr_block = 0;
    assign fifo_intf_616.finish = finish;
    csv_file_dump fifo_csv_dumper_616;
    csv_file_dump cstatus_csv_dumper_616;
    df_fifo_monitor fifo_monitor_616;
    df_fifo_intf fifo_intf_617(clock,reset);
    assign fifo_intf_617.rd_en = AESL_inst_myproject.layer2_out_616_U.if_read & AESL_inst_myproject.layer2_out_616_U.if_empty_n;
    assign fifo_intf_617.wr_en = AESL_inst_myproject.layer2_out_616_U.if_write & AESL_inst_myproject.layer2_out_616_U.if_full_n;
    assign fifo_intf_617.fifo_rd_block = 0;
    assign fifo_intf_617.fifo_wr_block = 0;
    assign fifo_intf_617.finish = finish;
    csv_file_dump fifo_csv_dumper_617;
    csv_file_dump cstatus_csv_dumper_617;
    df_fifo_monitor fifo_monitor_617;
    df_fifo_intf fifo_intf_618(clock,reset);
    assign fifo_intf_618.rd_en = AESL_inst_myproject.layer2_out_617_U.if_read & AESL_inst_myproject.layer2_out_617_U.if_empty_n;
    assign fifo_intf_618.wr_en = AESL_inst_myproject.layer2_out_617_U.if_write & AESL_inst_myproject.layer2_out_617_U.if_full_n;
    assign fifo_intf_618.fifo_rd_block = 0;
    assign fifo_intf_618.fifo_wr_block = 0;
    assign fifo_intf_618.finish = finish;
    csv_file_dump fifo_csv_dumper_618;
    csv_file_dump cstatus_csv_dumper_618;
    df_fifo_monitor fifo_monitor_618;
    df_fifo_intf fifo_intf_619(clock,reset);
    assign fifo_intf_619.rd_en = AESL_inst_myproject.layer2_out_618_U.if_read & AESL_inst_myproject.layer2_out_618_U.if_empty_n;
    assign fifo_intf_619.wr_en = AESL_inst_myproject.layer2_out_618_U.if_write & AESL_inst_myproject.layer2_out_618_U.if_full_n;
    assign fifo_intf_619.fifo_rd_block = 0;
    assign fifo_intf_619.fifo_wr_block = 0;
    assign fifo_intf_619.finish = finish;
    csv_file_dump fifo_csv_dumper_619;
    csv_file_dump cstatus_csv_dumper_619;
    df_fifo_monitor fifo_monitor_619;
    df_fifo_intf fifo_intf_620(clock,reset);
    assign fifo_intf_620.rd_en = AESL_inst_myproject.layer2_out_619_U.if_read & AESL_inst_myproject.layer2_out_619_U.if_empty_n;
    assign fifo_intf_620.wr_en = AESL_inst_myproject.layer2_out_619_U.if_write & AESL_inst_myproject.layer2_out_619_U.if_full_n;
    assign fifo_intf_620.fifo_rd_block = 0;
    assign fifo_intf_620.fifo_wr_block = 0;
    assign fifo_intf_620.finish = finish;
    csv_file_dump fifo_csv_dumper_620;
    csv_file_dump cstatus_csv_dumper_620;
    df_fifo_monitor fifo_monitor_620;
    df_fifo_intf fifo_intf_621(clock,reset);
    assign fifo_intf_621.rd_en = AESL_inst_myproject.layer2_out_620_U.if_read & AESL_inst_myproject.layer2_out_620_U.if_empty_n;
    assign fifo_intf_621.wr_en = AESL_inst_myproject.layer2_out_620_U.if_write & AESL_inst_myproject.layer2_out_620_U.if_full_n;
    assign fifo_intf_621.fifo_rd_block = 0;
    assign fifo_intf_621.fifo_wr_block = 0;
    assign fifo_intf_621.finish = finish;
    csv_file_dump fifo_csv_dumper_621;
    csv_file_dump cstatus_csv_dumper_621;
    df_fifo_monitor fifo_monitor_621;
    df_fifo_intf fifo_intf_622(clock,reset);
    assign fifo_intf_622.rd_en = AESL_inst_myproject.layer2_out_621_U.if_read & AESL_inst_myproject.layer2_out_621_U.if_empty_n;
    assign fifo_intf_622.wr_en = AESL_inst_myproject.layer2_out_621_U.if_write & AESL_inst_myproject.layer2_out_621_U.if_full_n;
    assign fifo_intf_622.fifo_rd_block = 0;
    assign fifo_intf_622.fifo_wr_block = 0;
    assign fifo_intf_622.finish = finish;
    csv_file_dump fifo_csv_dumper_622;
    csv_file_dump cstatus_csv_dumper_622;
    df_fifo_monitor fifo_monitor_622;
    df_fifo_intf fifo_intf_623(clock,reset);
    assign fifo_intf_623.rd_en = AESL_inst_myproject.layer2_out_622_U.if_read & AESL_inst_myproject.layer2_out_622_U.if_empty_n;
    assign fifo_intf_623.wr_en = AESL_inst_myproject.layer2_out_622_U.if_write & AESL_inst_myproject.layer2_out_622_U.if_full_n;
    assign fifo_intf_623.fifo_rd_block = 0;
    assign fifo_intf_623.fifo_wr_block = 0;
    assign fifo_intf_623.finish = finish;
    csv_file_dump fifo_csv_dumper_623;
    csv_file_dump cstatus_csv_dumper_623;
    df_fifo_monitor fifo_monitor_623;
    df_fifo_intf fifo_intf_624(clock,reset);
    assign fifo_intf_624.rd_en = AESL_inst_myproject.layer2_out_623_U.if_read & AESL_inst_myproject.layer2_out_623_U.if_empty_n;
    assign fifo_intf_624.wr_en = AESL_inst_myproject.layer2_out_623_U.if_write & AESL_inst_myproject.layer2_out_623_U.if_full_n;
    assign fifo_intf_624.fifo_rd_block = 0;
    assign fifo_intf_624.fifo_wr_block = 0;
    assign fifo_intf_624.finish = finish;
    csv_file_dump fifo_csv_dumper_624;
    csv_file_dump cstatus_csv_dumper_624;
    df_fifo_monitor fifo_monitor_624;
    df_fifo_intf fifo_intf_625(clock,reset);
    assign fifo_intf_625.rd_en = AESL_inst_myproject.layer2_out_624_U.if_read & AESL_inst_myproject.layer2_out_624_U.if_empty_n;
    assign fifo_intf_625.wr_en = AESL_inst_myproject.layer2_out_624_U.if_write & AESL_inst_myproject.layer2_out_624_U.if_full_n;
    assign fifo_intf_625.fifo_rd_block = 0;
    assign fifo_intf_625.fifo_wr_block = 0;
    assign fifo_intf_625.finish = finish;
    csv_file_dump fifo_csv_dumper_625;
    csv_file_dump cstatus_csv_dumper_625;
    df_fifo_monitor fifo_monitor_625;
    df_fifo_intf fifo_intf_626(clock,reset);
    assign fifo_intf_626.rd_en = AESL_inst_myproject.layer2_out_625_U.if_read & AESL_inst_myproject.layer2_out_625_U.if_empty_n;
    assign fifo_intf_626.wr_en = AESL_inst_myproject.layer2_out_625_U.if_write & AESL_inst_myproject.layer2_out_625_U.if_full_n;
    assign fifo_intf_626.fifo_rd_block = 0;
    assign fifo_intf_626.fifo_wr_block = 0;
    assign fifo_intf_626.finish = finish;
    csv_file_dump fifo_csv_dumper_626;
    csv_file_dump cstatus_csv_dumper_626;
    df_fifo_monitor fifo_monitor_626;
    df_fifo_intf fifo_intf_627(clock,reset);
    assign fifo_intf_627.rd_en = AESL_inst_myproject.layer2_out_626_U.if_read & AESL_inst_myproject.layer2_out_626_U.if_empty_n;
    assign fifo_intf_627.wr_en = AESL_inst_myproject.layer2_out_626_U.if_write & AESL_inst_myproject.layer2_out_626_U.if_full_n;
    assign fifo_intf_627.fifo_rd_block = 0;
    assign fifo_intf_627.fifo_wr_block = 0;
    assign fifo_intf_627.finish = finish;
    csv_file_dump fifo_csv_dumper_627;
    csv_file_dump cstatus_csv_dumper_627;
    df_fifo_monitor fifo_monitor_627;
    df_fifo_intf fifo_intf_628(clock,reset);
    assign fifo_intf_628.rd_en = AESL_inst_myproject.layer2_out_627_U.if_read & AESL_inst_myproject.layer2_out_627_U.if_empty_n;
    assign fifo_intf_628.wr_en = AESL_inst_myproject.layer2_out_627_U.if_write & AESL_inst_myproject.layer2_out_627_U.if_full_n;
    assign fifo_intf_628.fifo_rd_block = 0;
    assign fifo_intf_628.fifo_wr_block = 0;
    assign fifo_intf_628.finish = finish;
    csv_file_dump fifo_csv_dumper_628;
    csv_file_dump cstatus_csv_dumper_628;
    df_fifo_monitor fifo_monitor_628;
    df_fifo_intf fifo_intf_629(clock,reset);
    assign fifo_intf_629.rd_en = AESL_inst_myproject.layer2_out_628_U.if_read & AESL_inst_myproject.layer2_out_628_U.if_empty_n;
    assign fifo_intf_629.wr_en = AESL_inst_myproject.layer2_out_628_U.if_write & AESL_inst_myproject.layer2_out_628_U.if_full_n;
    assign fifo_intf_629.fifo_rd_block = 0;
    assign fifo_intf_629.fifo_wr_block = 0;
    assign fifo_intf_629.finish = finish;
    csv_file_dump fifo_csv_dumper_629;
    csv_file_dump cstatus_csv_dumper_629;
    df_fifo_monitor fifo_monitor_629;
    df_fifo_intf fifo_intf_630(clock,reset);
    assign fifo_intf_630.rd_en = AESL_inst_myproject.layer2_out_629_U.if_read & AESL_inst_myproject.layer2_out_629_U.if_empty_n;
    assign fifo_intf_630.wr_en = AESL_inst_myproject.layer2_out_629_U.if_write & AESL_inst_myproject.layer2_out_629_U.if_full_n;
    assign fifo_intf_630.fifo_rd_block = 0;
    assign fifo_intf_630.fifo_wr_block = 0;
    assign fifo_intf_630.finish = finish;
    csv_file_dump fifo_csv_dumper_630;
    csv_file_dump cstatus_csv_dumper_630;
    df_fifo_monitor fifo_monitor_630;
    df_fifo_intf fifo_intf_631(clock,reset);
    assign fifo_intf_631.rd_en = AESL_inst_myproject.layer2_out_630_U.if_read & AESL_inst_myproject.layer2_out_630_U.if_empty_n;
    assign fifo_intf_631.wr_en = AESL_inst_myproject.layer2_out_630_U.if_write & AESL_inst_myproject.layer2_out_630_U.if_full_n;
    assign fifo_intf_631.fifo_rd_block = 0;
    assign fifo_intf_631.fifo_wr_block = 0;
    assign fifo_intf_631.finish = finish;
    csv_file_dump fifo_csv_dumper_631;
    csv_file_dump cstatus_csv_dumper_631;
    df_fifo_monitor fifo_monitor_631;
    df_fifo_intf fifo_intf_632(clock,reset);
    assign fifo_intf_632.rd_en = AESL_inst_myproject.layer2_out_631_U.if_read & AESL_inst_myproject.layer2_out_631_U.if_empty_n;
    assign fifo_intf_632.wr_en = AESL_inst_myproject.layer2_out_631_U.if_write & AESL_inst_myproject.layer2_out_631_U.if_full_n;
    assign fifo_intf_632.fifo_rd_block = 0;
    assign fifo_intf_632.fifo_wr_block = 0;
    assign fifo_intf_632.finish = finish;
    csv_file_dump fifo_csv_dumper_632;
    csv_file_dump cstatus_csv_dumper_632;
    df_fifo_monitor fifo_monitor_632;
    df_fifo_intf fifo_intf_633(clock,reset);
    assign fifo_intf_633.rd_en = AESL_inst_myproject.layer2_out_632_U.if_read & AESL_inst_myproject.layer2_out_632_U.if_empty_n;
    assign fifo_intf_633.wr_en = AESL_inst_myproject.layer2_out_632_U.if_write & AESL_inst_myproject.layer2_out_632_U.if_full_n;
    assign fifo_intf_633.fifo_rd_block = 0;
    assign fifo_intf_633.fifo_wr_block = 0;
    assign fifo_intf_633.finish = finish;
    csv_file_dump fifo_csv_dumper_633;
    csv_file_dump cstatus_csv_dumper_633;
    df_fifo_monitor fifo_monitor_633;
    df_fifo_intf fifo_intf_634(clock,reset);
    assign fifo_intf_634.rd_en = AESL_inst_myproject.layer2_out_633_U.if_read & AESL_inst_myproject.layer2_out_633_U.if_empty_n;
    assign fifo_intf_634.wr_en = AESL_inst_myproject.layer2_out_633_U.if_write & AESL_inst_myproject.layer2_out_633_U.if_full_n;
    assign fifo_intf_634.fifo_rd_block = 0;
    assign fifo_intf_634.fifo_wr_block = 0;
    assign fifo_intf_634.finish = finish;
    csv_file_dump fifo_csv_dumper_634;
    csv_file_dump cstatus_csv_dumper_634;
    df_fifo_monitor fifo_monitor_634;
    df_fifo_intf fifo_intf_635(clock,reset);
    assign fifo_intf_635.rd_en = AESL_inst_myproject.layer2_out_634_U.if_read & AESL_inst_myproject.layer2_out_634_U.if_empty_n;
    assign fifo_intf_635.wr_en = AESL_inst_myproject.layer2_out_634_U.if_write & AESL_inst_myproject.layer2_out_634_U.if_full_n;
    assign fifo_intf_635.fifo_rd_block = 0;
    assign fifo_intf_635.fifo_wr_block = 0;
    assign fifo_intf_635.finish = finish;
    csv_file_dump fifo_csv_dumper_635;
    csv_file_dump cstatus_csv_dumper_635;
    df_fifo_monitor fifo_monitor_635;
    df_fifo_intf fifo_intf_636(clock,reset);
    assign fifo_intf_636.rd_en = AESL_inst_myproject.layer2_out_635_U.if_read & AESL_inst_myproject.layer2_out_635_U.if_empty_n;
    assign fifo_intf_636.wr_en = AESL_inst_myproject.layer2_out_635_U.if_write & AESL_inst_myproject.layer2_out_635_U.if_full_n;
    assign fifo_intf_636.fifo_rd_block = 0;
    assign fifo_intf_636.fifo_wr_block = 0;
    assign fifo_intf_636.finish = finish;
    csv_file_dump fifo_csv_dumper_636;
    csv_file_dump cstatus_csv_dumper_636;
    df_fifo_monitor fifo_monitor_636;
    df_fifo_intf fifo_intf_637(clock,reset);
    assign fifo_intf_637.rd_en = AESL_inst_myproject.layer2_out_636_U.if_read & AESL_inst_myproject.layer2_out_636_U.if_empty_n;
    assign fifo_intf_637.wr_en = AESL_inst_myproject.layer2_out_636_U.if_write & AESL_inst_myproject.layer2_out_636_U.if_full_n;
    assign fifo_intf_637.fifo_rd_block = 0;
    assign fifo_intf_637.fifo_wr_block = 0;
    assign fifo_intf_637.finish = finish;
    csv_file_dump fifo_csv_dumper_637;
    csv_file_dump cstatus_csv_dumper_637;
    df_fifo_monitor fifo_monitor_637;
    df_fifo_intf fifo_intf_638(clock,reset);
    assign fifo_intf_638.rd_en = AESL_inst_myproject.layer2_out_637_U.if_read & AESL_inst_myproject.layer2_out_637_U.if_empty_n;
    assign fifo_intf_638.wr_en = AESL_inst_myproject.layer2_out_637_U.if_write & AESL_inst_myproject.layer2_out_637_U.if_full_n;
    assign fifo_intf_638.fifo_rd_block = 0;
    assign fifo_intf_638.fifo_wr_block = 0;
    assign fifo_intf_638.finish = finish;
    csv_file_dump fifo_csv_dumper_638;
    csv_file_dump cstatus_csv_dumper_638;
    df_fifo_monitor fifo_monitor_638;
    df_fifo_intf fifo_intf_639(clock,reset);
    assign fifo_intf_639.rd_en = AESL_inst_myproject.layer2_out_638_U.if_read & AESL_inst_myproject.layer2_out_638_U.if_empty_n;
    assign fifo_intf_639.wr_en = AESL_inst_myproject.layer2_out_638_U.if_write & AESL_inst_myproject.layer2_out_638_U.if_full_n;
    assign fifo_intf_639.fifo_rd_block = 0;
    assign fifo_intf_639.fifo_wr_block = 0;
    assign fifo_intf_639.finish = finish;
    csv_file_dump fifo_csv_dumper_639;
    csv_file_dump cstatus_csv_dumper_639;
    df_fifo_monitor fifo_monitor_639;
    df_fifo_intf fifo_intf_640(clock,reset);
    assign fifo_intf_640.rd_en = AESL_inst_myproject.layer2_out_639_U.if_read & AESL_inst_myproject.layer2_out_639_U.if_empty_n;
    assign fifo_intf_640.wr_en = AESL_inst_myproject.layer2_out_639_U.if_write & AESL_inst_myproject.layer2_out_639_U.if_full_n;
    assign fifo_intf_640.fifo_rd_block = 0;
    assign fifo_intf_640.fifo_wr_block = 0;
    assign fifo_intf_640.finish = finish;
    csv_file_dump fifo_csv_dumper_640;
    csv_file_dump cstatus_csv_dumper_640;
    df_fifo_monitor fifo_monitor_640;
    df_fifo_intf fifo_intf_641(clock,reset);
    assign fifo_intf_641.rd_en = AESL_inst_myproject.layer2_out_640_U.if_read & AESL_inst_myproject.layer2_out_640_U.if_empty_n;
    assign fifo_intf_641.wr_en = AESL_inst_myproject.layer2_out_640_U.if_write & AESL_inst_myproject.layer2_out_640_U.if_full_n;
    assign fifo_intf_641.fifo_rd_block = 0;
    assign fifo_intf_641.fifo_wr_block = 0;
    assign fifo_intf_641.finish = finish;
    csv_file_dump fifo_csv_dumper_641;
    csv_file_dump cstatus_csv_dumper_641;
    df_fifo_monitor fifo_monitor_641;
    df_fifo_intf fifo_intf_642(clock,reset);
    assign fifo_intf_642.rd_en = AESL_inst_myproject.layer2_out_641_U.if_read & AESL_inst_myproject.layer2_out_641_U.if_empty_n;
    assign fifo_intf_642.wr_en = AESL_inst_myproject.layer2_out_641_U.if_write & AESL_inst_myproject.layer2_out_641_U.if_full_n;
    assign fifo_intf_642.fifo_rd_block = 0;
    assign fifo_intf_642.fifo_wr_block = 0;
    assign fifo_intf_642.finish = finish;
    csv_file_dump fifo_csv_dumper_642;
    csv_file_dump cstatus_csv_dumper_642;
    df_fifo_monitor fifo_monitor_642;
    df_fifo_intf fifo_intf_643(clock,reset);
    assign fifo_intf_643.rd_en = AESL_inst_myproject.layer2_out_642_U.if_read & AESL_inst_myproject.layer2_out_642_U.if_empty_n;
    assign fifo_intf_643.wr_en = AESL_inst_myproject.layer2_out_642_U.if_write & AESL_inst_myproject.layer2_out_642_U.if_full_n;
    assign fifo_intf_643.fifo_rd_block = 0;
    assign fifo_intf_643.fifo_wr_block = 0;
    assign fifo_intf_643.finish = finish;
    csv_file_dump fifo_csv_dumper_643;
    csv_file_dump cstatus_csv_dumper_643;
    df_fifo_monitor fifo_monitor_643;
    df_fifo_intf fifo_intf_644(clock,reset);
    assign fifo_intf_644.rd_en = AESL_inst_myproject.layer2_out_643_U.if_read & AESL_inst_myproject.layer2_out_643_U.if_empty_n;
    assign fifo_intf_644.wr_en = AESL_inst_myproject.layer2_out_643_U.if_write & AESL_inst_myproject.layer2_out_643_U.if_full_n;
    assign fifo_intf_644.fifo_rd_block = 0;
    assign fifo_intf_644.fifo_wr_block = 0;
    assign fifo_intf_644.finish = finish;
    csv_file_dump fifo_csv_dumper_644;
    csv_file_dump cstatus_csv_dumper_644;
    df_fifo_monitor fifo_monitor_644;
    df_fifo_intf fifo_intf_645(clock,reset);
    assign fifo_intf_645.rd_en = AESL_inst_myproject.layer2_out_644_U.if_read & AESL_inst_myproject.layer2_out_644_U.if_empty_n;
    assign fifo_intf_645.wr_en = AESL_inst_myproject.layer2_out_644_U.if_write & AESL_inst_myproject.layer2_out_644_U.if_full_n;
    assign fifo_intf_645.fifo_rd_block = 0;
    assign fifo_intf_645.fifo_wr_block = 0;
    assign fifo_intf_645.finish = finish;
    csv_file_dump fifo_csv_dumper_645;
    csv_file_dump cstatus_csv_dumper_645;
    df_fifo_monitor fifo_monitor_645;
    df_fifo_intf fifo_intf_646(clock,reset);
    assign fifo_intf_646.rd_en = AESL_inst_myproject.layer2_out_645_U.if_read & AESL_inst_myproject.layer2_out_645_U.if_empty_n;
    assign fifo_intf_646.wr_en = AESL_inst_myproject.layer2_out_645_U.if_write & AESL_inst_myproject.layer2_out_645_U.if_full_n;
    assign fifo_intf_646.fifo_rd_block = 0;
    assign fifo_intf_646.fifo_wr_block = 0;
    assign fifo_intf_646.finish = finish;
    csv_file_dump fifo_csv_dumper_646;
    csv_file_dump cstatus_csv_dumper_646;
    df_fifo_monitor fifo_monitor_646;
    df_fifo_intf fifo_intf_647(clock,reset);
    assign fifo_intf_647.rd_en = AESL_inst_myproject.layer2_out_646_U.if_read & AESL_inst_myproject.layer2_out_646_U.if_empty_n;
    assign fifo_intf_647.wr_en = AESL_inst_myproject.layer2_out_646_U.if_write & AESL_inst_myproject.layer2_out_646_U.if_full_n;
    assign fifo_intf_647.fifo_rd_block = 0;
    assign fifo_intf_647.fifo_wr_block = 0;
    assign fifo_intf_647.finish = finish;
    csv_file_dump fifo_csv_dumper_647;
    csv_file_dump cstatus_csv_dumper_647;
    df_fifo_monitor fifo_monitor_647;
    df_fifo_intf fifo_intf_648(clock,reset);
    assign fifo_intf_648.rd_en = AESL_inst_myproject.layer2_out_647_U.if_read & AESL_inst_myproject.layer2_out_647_U.if_empty_n;
    assign fifo_intf_648.wr_en = AESL_inst_myproject.layer2_out_647_U.if_write & AESL_inst_myproject.layer2_out_647_U.if_full_n;
    assign fifo_intf_648.fifo_rd_block = 0;
    assign fifo_intf_648.fifo_wr_block = 0;
    assign fifo_intf_648.finish = finish;
    csv_file_dump fifo_csv_dumper_648;
    csv_file_dump cstatus_csv_dumper_648;
    df_fifo_monitor fifo_monitor_648;
    df_fifo_intf fifo_intf_649(clock,reset);
    assign fifo_intf_649.rd_en = AESL_inst_myproject.layer2_out_648_U.if_read & AESL_inst_myproject.layer2_out_648_U.if_empty_n;
    assign fifo_intf_649.wr_en = AESL_inst_myproject.layer2_out_648_U.if_write & AESL_inst_myproject.layer2_out_648_U.if_full_n;
    assign fifo_intf_649.fifo_rd_block = 0;
    assign fifo_intf_649.fifo_wr_block = 0;
    assign fifo_intf_649.finish = finish;
    csv_file_dump fifo_csv_dumper_649;
    csv_file_dump cstatus_csv_dumper_649;
    df_fifo_monitor fifo_monitor_649;
    df_fifo_intf fifo_intf_650(clock,reset);
    assign fifo_intf_650.rd_en = AESL_inst_myproject.layer2_out_649_U.if_read & AESL_inst_myproject.layer2_out_649_U.if_empty_n;
    assign fifo_intf_650.wr_en = AESL_inst_myproject.layer2_out_649_U.if_write & AESL_inst_myproject.layer2_out_649_U.if_full_n;
    assign fifo_intf_650.fifo_rd_block = 0;
    assign fifo_intf_650.fifo_wr_block = 0;
    assign fifo_intf_650.finish = finish;
    csv_file_dump fifo_csv_dumper_650;
    csv_file_dump cstatus_csv_dumper_650;
    df_fifo_monitor fifo_monitor_650;
    df_fifo_intf fifo_intf_651(clock,reset);
    assign fifo_intf_651.rd_en = AESL_inst_myproject.layer2_out_650_U.if_read & AESL_inst_myproject.layer2_out_650_U.if_empty_n;
    assign fifo_intf_651.wr_en = AESL_inst_myproject.layer2_out_650_U.if_write & AESL_inst_myproject.layer2_out_650_U.if_full_n;
    assign fifo_intf_651.fifo_rd_block = 0;
    assign fifo_intf_651.fifo_wr_block = 0;
    assign fifo_intf_651.finish = finish;
    csv_file_dump fifo_csv_dumper_651;
    csv_file_dump cstatus_csv_dumper_651;
    df_fifo_monitor fifo_monitor_651;
    df_fifo_intf fifo_intf_652(clock,reset);
    assign fifo_intf_652.rd_en = AESL_inst_myproject.layer2_out_651_U.if_read & AESL_inst_myproject.layer2_out_651_U.if_empty_n;
    assign fifo_intf_652.wr_en = AESL_inst_myproject.layer2_out_651_U.if_write & AESL_inst_myproject.layer2_out_651_U.if_full_n;
    assign fifo_intf_652.fifo_rd_block = 0;
    assign fifo_intf_652.fifo_wr_block = 0;
    assign fifo_intf_652.finish = finish;
    csv_file_dump fifo_csv_dumper_652;
    csv_file_dump cstatus_csv_dumper_652;
    df_fifo_monitor fifo_monitor_652;
    df_fifo_intf fifo_intf_653(clock,reset);
    assign fifo_intf_653.rd_en = AESL_inst_myproject.layer2_out_652_U.if_read & AESL_inst_myproject.layer2_out_652_U.if_empty_n;
    assign fifo_intf_653.wr_en = AESL_inst_myproject.layer2_out_652_U.if_write & AESL_inst_myproject.layer2_out_652_U.if_full_n;
    assign fifo_intf_653.fifo_rd_block = 0;
    assign fifo_intf_653.fifo_wr_block = 0;
    assign fifo_intf_653.finish = finish;
    csv_file_dump fifo_csv_dumper_653;
    csv_file_dump cstatus_csv_dumper_653;
    df_fifo_monitor fifo_monitor_653;
    df_fifo_intf fifo_intf_654(clock,reset);
    assign fifo_intf_654.rd_en = AESL_inst_myproject.layer2_out_653_U.if_read & AESL_inst_myproject.layer2_out_653_U.if_empty_n;
    assign fifo_intf_654.wr_en = AESL_inst_myproject.layer2_out_653_U.if_write & AESL_inst_myproject.layer2_out_653_U.if_full_n;
    assign fifo_intf_654.fifo_rd_block = 0;
    assign fifo_intf_654.fifo_wr_block = 0;
    assign fifo_intf_654.finish = finish;
    csv_file_dump fifo_csv_dumper_654;
    csv_file_dump cstatus_csv_dumper_654;
    df_fifo_monitor fifo_monitor_654;
    df_fifo_intf fifo_intf_655(clock,reset);
    assign fifo_intf_655.rd_en = AESL_inst_myproject.layer2_out_654_U.if_read & AESL_inst_myproject.layer2_out_654_U.if_empty_n;
    assign fifo_intf_655.wr_en = AESL_inst_myproject.layer2_out_654_U.if_write & AESL_inst_myproject.layer2_out_654_U.if_full_n;
    assign fifo_intf_655.fifo_rd_block = 0;
    assign fifo_intf_655.fifo_wr_block = 0;
    assign fifo_intf_655.finish = finish;
    csv_file_dump fifo_csv_dumper_655;
    csv_file_dump cstatus_csv_dumper_655;
    df_fifo_monitor fifo_monitor_655;
    df_fifo_intf fifo_intf_656(clock,reset);
    assign fifo_intf_656.rd_en = AESL_inst_myproject.layer2_out_655_U.if_read & AESL_inst_myproject.layer2_out_655_U.if_empty_n;
    assign fifo_intf_656.wr_en = AESL_inst_myproject.layer2_out_655_U.if_write & AESL_inst_myproject.layer2_out_655_U.if_full_n;
    assign fifo_intf_656.fifo_rd_block = 0;
    assign fifo_intf_656.fifo_wr_block = 0;
    assign fifo_intf_656.finish = finish;
    csv_file_dump fifo_csv_dumper_656;
    csv_file_dump cstatus_csv_dumper_656;
    df_fifo_monitor fifo_monitor_656;
    df_fifo_intf fifo_intf_657(clock,reset);
    assign fifo_intf_657.rd_en = AESL_inst_myproject.layer2_out_656_U.if_read & AESL_inst_myproject.layer2_out_656_U.if_empty_n;
    assign fifo_intf_657.wr_en = AESL_inst_myproject.layer2_out_656_U.if_write & AESL_inst_myproject.layer2_out_656_U.if_full_n;
    assign fifo_intf_657.fifo_rd_block = 0;
    assign fifo_intf_657.fifo_wr_block = 0;
    assign fifo_intf_657.finish = finish;
    csv_file_dump fifo_csv_dumper_657;
    csv_file_dump cstatus_csv_dumper_657;
    df_fifo_monitor fifo_monitor_657;
    df_fifo_intf fifo_intf_658(clock,reset);
    assign fifo_intf_658.rd_en = AESL_inst_myproject.layer2_out_657_U.if_read & AESL_inst_myproject.layer2_out_657_U.if_empty_n;
    assign fifo_intf_658.wr_en = AESL_inst_myproject.layer2_out_657_U.if_write & AESL_inst_myproject.layer2_out_657_U.if_full_n;
    assign fifo_intf_658.fifo_rd_block = 0;
    assign fifo_intf_658.fifo_wr_block = 0;
    assign fifo_intf_658.finish = finish;
    csv_file_dump fifo_csv_dumper_658;
    csv_file_dump cstatus_csv_dumper_658;
    df_fifo_monitor fifo_monitor_658;
    df_fifo_intf fifo_intf_659(clock,reset);
    assign fifo_intf_659.rd_en = AESL_inst_myproject.layer2_out_658_U.if_read & AESL_inst_myproject.layer2_out_658_U.if_empty_n;
    assign fifo_intf_659.wr_en = AESL_inst_myproject.layer2_out_658_U.if_write & AESL_inst_myproject.layer2_out_658_U.if_full_n;
    assign fifo_intf_659.fifo_rd_block = 0;
    assign fifo_intf_659.fifo_wr_block = 0;
    assign fifo_intf_659.finish = finish;
    csv_file_dump fifo_csv_dumper_659;
    csv_file_dump cstatus_csv_dumper_659;
    df_fifo_monitor fifo_monitor_659;
    df_fifo_intf fifo_intf_660(clock,reset);
    assign fifo_intf_660.rd_en = AESL_inst_myproject.layer2_out_659_U.if_read & AESL_inst_myproject.layer2_out_659_U.if_empty_n;
    assign fifo_intf_660.wr_en = AESL_inst_myproject.layer2_out_659_U.if_write & AESL_inst_myproject.layer2_out_659_U.if_full_n;
    assign fifo_intf_660.fifo_rd_block = 0;
    assign fifo_intf_660.fifo_wr_block = 0;
    assign fifo_intf_660.finish = finish;
    csv_file_dump fifo_csv_dumper_660;
    csv_file_dump cstatus_csv_dumper_660;
    df_fifo_monitor fifo_monitor_660;
    df_fifo_intf fifo_intf_661(clock,reset);
    assign fifo_intf_661.rd_en = AESL_inst_myproject.layer2_out_660_U.if_read & AESL_inst_myproject.layer2_out_660_U.if_empty_n;
    assign fifo_intf_661.wr_en = AESL_inst_myproject.layer2_out_660_U.if_write & AESL_inst_myproject.layer2_out_660_U.if_full_n;
    assign fifo_intf_661.fifo_rd_block = 0;
    assign fifo_intf_661.fifo_wr_block = 0;
    assign fifo_intf_661.finish = finish;
    csv_file_dump fifo_csv_dumper_661;
    csv_file_dump cstatus_csv_dumper_661;
    df_fifo_monitor fifo_monitor_661;
    df_fifo_intf fifo_intf_662(clock,reset);
    assign fifo_intf_662.rd_en = AESL_inst_myproject.layer2_out_661_U.if_read & AESL_inst_myproject.layer2_out_661_U.if_empty_n;
    assign fifo_intf_662.wr_en = AESL_inst_myproject.layer2_out_661_U.if_write & AESL_inst_myproject.layer2_out_661_U.if_full_n;
    assign fifo_intf_662.fifo_rd_block = 0;
    assign fifo_intf_662.fifo_wr_block = 0;
    assign fifo_intf_662.finish = finish;
    csv_file_dump fifo_csv_dumper_662;
    csv_file_dump cstatus_csv_dumper_662;
    df_fifo_monitor fifo_monitor_662;
    df_fifo_intf fifo_intf_663(clock,reset);
    assign fifo_intf_663.rd_en = AESL_inst_myproject.layer2_out_662_U.if_read & AESL_inst_myproject.layer2_out_662_U.if_empty_n;
    assign fifo_intf_663.wr_en = AESL_inst_myproject.layer2_out_662_U.if_write & AESL_inst_myproject.layer2_out_662_U.if_full_n;
    assign fifo_intf_663.fifo_rd_block = 0;
    assign fifo_intf_663.fifo_wr_block = 0;
    assign fifo_intf_663.finish = finish;
    csv_file_dump fifo_csv_dumper_663;
    csv_file_dump cstatus_csv_dumper_663;
    df_fifo_monitor fifo_monitor_663;
    df_fifo_intf fifo_intf_664(clock,reset);
    assign fifo_intf_664.rd_en = AESL_inst_myproject.layer2_out_663_U.if_read & AESL_inst_myproject.layer2_out_663_U.if_empty_n;
    assign fifo_intf_664.wr_en = AESL_inst_myproject.layer2_out_663_U.if_write & AESL_inst_myproject.layer2_out_663_U.if_full_n;
    assign fifo_intf_664.fifo_rd_block = 0;
    assign fifo_intf_664.fifo_wr_block = 0;
    assign fifo_intf_664.finish = finish;
    csv_file_dump fifo_csv_dumper_664;
    csv_file_dump cstatus_csv_dumper_664;
    df_fifo_monitor fifo_monitor_664;
    df_fifo_intf fifo_intf_665(clock,reset);
    assign fifo_intf_665.rd_en = AESL_inst_myproject.layer2_out_664_U.if_read & AESL_inst_myproject.layer2_out_664_U.if_empty_n;
    assign fifo_intf_665.wr_en = AESL_inst_myproject.layer2_out_664_U.if_write & AESL_inst_myproject.layer2_out_664_U.if_full_n;
    assign fifo_intf_665.fifo_rd_block = 0;
    assign fifo_intf_665.fifo_wr_block = 0;
    assign fifo_intf_665.finish = finish;
    csv_file_dump fifo_csv_dumper_665;
    csv_file_dump cstatus_csv_dumper_665;
    df_fifo_monitor fifo_monitor_665;
    df_fifo_intf fifo_intf_666(clock,reset);
    assign fifo_intf_666.rd_en = AESL_inst_myproject.layer2_out_665_U.if_read & AESL_inst_myproject.layer2_out_665_U.if_empty_n;
    assign fifo_intf_666.wr_en = AESL_inst_myproject.layer2_out_665_U.if_write & AESL_inst_myproject.layer2_out_665_U.if_full_n;
    assign fifo_intf_666.fifo_rd_block = 0;
    assign fifo_intf_666.fifo_wr_block = 0;
    assign fifo_intf_666.finish = finish;
    csv_file_dump fifo_csv_dumper_666;
    csv_file_dump cstatus_csv_dumper_666;
    df_fifo_monitor fifo_monitor_666;
    df_fifo_intf fifo_intf_667(clock,reset);
    assign fifo_intf_667.rd_en = AESL_inst_myproject.layer2_out_666_U.if_read & AESL_inst_myproject.layer2_out_666_U.if_empty_n;
    assign fifo_intf_667.wr_en = AESL_inst_myproject.layer2_out_666_U.if_write & AESL_inst_myproject.layer2_out_666_U.if_full_n;
    assign fifo_intf_667.fifo_rd_block = 0;
    assign fifo_intf_667.fifo_wr_block = 0;
    assign fifo_intf_667.finish = finish;
    csv_file_dump fifo_csv_dumper_667;
    csv_file_dump cstatus_csv_dumper_667;
    df_fifo_monitor fifo_monitor_667;
    df_fifo_intf fifo_intf_668(clock,reset);
    assign fifo_intf_668.rd_en = AESL_inst_myproject.layer2_out_667_U.if_read & AESL_inst_myproject.layer2_out_667_U.if_empty_n;
    assign fifo_intf_668.wr_en = AESL_inst_myproject.layer2_out_667_U.if_write & AESL_inst_myproject.layer2_out_667_U.if_full_n;
    assign fifo_intf_668.fifo_rd_block = 0;
    assign fifo_intf_668.fifo_wr_block = 0;
    assign fifo_intf_668.finish = finish;
    csv_file_dump fifo_csv_dumper_668;
    csv_file_dump cstatus_csv_dumper_668;
    df_fifo_monitor fifo_monitor_668;
    df_fifo_intf fifo_intf_669(clock,reset);
    assign fifo_intf_669.rd_en = AESL_inst_myproject.layer2_out_668_U.if_read & AESL_inst_myproject.layer2_out_668_U.if_empty_n;
    assign fifo_intf_669.wr_en = AESL_inst_myproject.layer2_out_668_U.if_write & AESL_inst_myproject.layer2_out_668_U.if_full_n;
    assign fifo_intf_669.fifo_rd_block = 0;
    assign fifo_intf_669.fifo_wr_block = 0;
    assign fifo_intf_669.finish = finish;
    csv_file_dump fifo_csv_dumper_669;
    csv_file_dump cstatus_csv_dumper_669;
    df_fifo_monitor fifo_monitor_669;
    df_fifo_intf fifo_intf_670(clock,reset);
    assign fifo_intf_670.rd_en = AESL_inst_myproject.layer2_out_669_U.if_read & AESL_inst_myproject.layer2_out_669_U.if_empty_n;
    assign fifo_intf_670.wr_en = AESL_inst_myproject.layer2_out_669_U.if_write & AESL_inst_myproject.layer2_out_669_U.if_full_n;
    assign fifo_intf_670.fifo_rd_block = 0;
    assign fifo_intf_670.fifo_wr_block = 0;
    assign fifo_intf_670.finish = finish;
    csv_file_dump fifo_csv_dumper_670;
    csv_file_dump cstatus_csv_dumper_670;
    df_fifo_monitor fifo_monitor_670;
    df_fifo_intf fifo_intf_671(clock,reset);
    assign fifo_intf_671.rd_en = AESL_inst_myproject.layer2_out_670_U.if_read & AESL_inst_myproject.layer2_out_670_U.if_empty_n;
    assign fifo_intf_671.wr_en = AESL_inst_myproject.layer2_out_670_U.if_write & AESL_inst_myproject.layer2_out_670_U.if_full_n;
    assign fifo_intf_671.fifo_rd_block = 0;
    assign fifo_intf_671.fifo_wr_block = 0;
    assign fifo_intf_671.finish = finish;
    csv_file_dump fifo_csv_dumper_671;
    csv_file_dump cstatus_csv_dumper_671;
    df_fifo_monitor fifo_monitor_671;
    df_fifo_intf fifo_intf_672(clock,reset);
    assign fifo_intf_672.rd_en = AESL_inst_myproject.layer2_out_671_U.if_read & AESL_inst_myproject.layer2_out_671_U.if_empty_n;
    assign fifo_intf_672.wr_en = AESL_inst_myproject.layer2_out_671_U.if_write & AESL_inst_myproject.layer2_out_671_U.if_full_n;
    assign fifo_intf_672.fifo_rd_block = 0;
    assign fifo_intf_672.fifo_wr_block = 0;
    assign fifo_intf_672.finish = finish;
    csv_file_dump fifo_csv_dumper_672;
    csv_file_dump cstatus_csv_dumper_672;
    df_fifo_monitor fifo_monitor_672;
    df_fifo_intf fifo_intf_673(clock,reset);
    assign fifo_intf_673.rd_en = AESL_inst_myproject.layer2_out_672_U.if_read & AESL_inst_myproject.layer2_out_672_U.if_empty_n;
    assign fifo_intf_673.wr_en = AESL_inst_myproject.layer2_out_672_U.if_write & AESL_inst_myproject.layer2_out_672_U.if_full_n;
    assign fifo_intf_673.fifo_rd_block = 0;
    assign fifo_intf_673.fifo_wr_block = 0;
    assign fifo_intf_673.finish = finish;
    csv_file_dump fifo_csv_dumper_673;
    csv_file_dump cstatus_csv_dumper_673;
    df_fifo_monitor fifo_monitor_673;
    df_fifo_intf fifo_intf_674(clock,reset);
    assign fifo_intf_674.rd_en = AESL_inst_myproject.layer2_out_673_U.if_read & AESL_inst_myproject.layer2_out_673_U.if_empty_n;
    assign fifo_intf_674.wr_en = AESL_inst_myproject.layer2_out_673_U.if_write & AESL_inst_myproject.layer2_out_673_U.if_full_n;
    assign fifo_intf_674.fifo_rd_block = 0;
    assign fifo_intf_674.fifo_wr_block = 0;
    assign fifo_intf_674.finish = finish;
    csv_file_dump fifo_csv_dumper_674;
    csv_file_dump cstatus_csv_dumper_674;
    df_fifo_monitor fifo_monitor_674;
    df_fifo_intf fifo_intf_675(clock,reset);
    assign fifo_intf_675.rd_en = AESL_inst_myproject.layer2_out_674_U.if_read & AESL_inst_myproject.layer2_out_674_U.if_empty_n;
    assign fifo_intf_675.wr_en = AESL_inst_myproject.layer2_out_674_U.if_write & AESL_inst_myproject.layer2_out_674_U.if_full_n;
    assign fifo_intf_675.fifo_rd_block = 0;
    assign fifo_intf_675.fifo_wr_block = 0;
    assign fifo_intf_675.finish = finish;
    csv_file_dump fifo_csv_dumper_675;
    csv_file_dump cstatus_csv_dumper_675;
    df_fifo_monitor fifo_monitor_675;
    df_fifo_intf fifo_intf_676(clock,reset);
    assign fifo_intf_676.rd_en = AESL_inst_myproject.layer2_out_675_U.if_read & AESL_inst_myproject.layer2_out_675_U.if_empty_n;
    assign fifo_intf_676.wr_en = AESL_inst_myproject.layer2_out_675_U.if_write & AESL_inst_myproject.layer2_out_675_U.if_full_n;
    assign fifo_intf_676.fifo_rd_block = 0;
    assign fifo_intf_676.fifo_wr_block = 0;
    assign fifo_intf_676.finish = finish;
    csv_file_dump fifo_csv_dumper_676;
    csv_file_dump cstatus_csv_dumper_676;
    df_fifo_monitor fifo_monitor_676;
    df_fifo_intf fifo_intf_677(clock,reset);
    assign fifo_intf_677.rd_en = AESL_inst_myproject.layer2_out_676_U.if_read & AESL_inst_myproject.layer2_out_676_U.if_empty_n;
    assign fifo_intf_677.wr_en = AESL_inst_myproject.layer2_out_676_U.if_write & AESL_inst_myproject.layer2_out_676_U.if_full_n;
    assign fifo_intf_677.fifo_rd_block = 0;
    assign fifo_intf_677.fifo_wr_block = 0;
    assign fifo_intf_677.finish = finish;
    csv_file_dump fifo_csv_dumper_677;
    csv_file_dump cstatus_csv_dumper_677;
    df_fifo_monitor fifo_monitor_677;
    df_fifo_intf fifo_intf_678(clock,reset);
    assign fifo_intf_678.rd_en = AESL_inst_myproject.layer2_out_677_U.if_read & AESL_inst_myproject.layer2_out_677_U.if_empty_n;
    assign fifo_intf_678.wr_en = AESL_inst_myproject.layer2_out_677_U.if_write & AESL_inst_myproject.layer2_out_677_U.if_full_n;
    assign fifo_intf_678.fifo_rd_block = 0;
    assign fifo_intf_678.fifo_wr_block = 0;
    assign fifo_intf_678.finish = finish;
    csv_file_dump fifo_csv_dumper_678;
    csv_file_dump cstatus_csv_dumper_678;
    df_fifo_monitor fifo_monitor_678;
    df_fifo_intf fifo_intf_679(clock,reset);
    assign fifo_intf_679.rd_en = AESL_inst_myproject.layer2_out_678_U.if_read & AESL_inst_myproject.layer2_out_678_U.if_empty_n;
    assign fifo_intf_679.wr_en = AESL_inst_myproject.layer2_out_678_U.if_write & AESL_inst_myproject.layer2_out_678_U.if_full_n;
    assign fifo_intf_679.fifo_rd_block = 0;
    assign fifo_intf_679.fifo_wr_block = 0;
    assign fifo_intf_679.finish = finish;
    csv_file_dump fifo_csv_dumper_679;
    csv_file_dump cstatus_csv_dumper_679;
    df_fifo_monitor fifo_monitor_679;
    df_fifo_intf fifo_intf_680(clock,reset);
    assign fifo_intf_680.rd_en = AESL_inst_myproject.layer2_out_679_U.if_read & AESL_inst_myproject.layer2_out_679_U.if_empty_n;
    assign fifo_intf_680.wr_en = AESL_inst_myproject.layer2_out_679_U.if_write & AESL_inst_myproject.layer2_out_679_U.if_full_n;
    assign fifo_intf_680.fifo_rd_block = 0;
    assign fifo_intf_680.fifo_wr_block = 0;
    assign fifo_intf_680.finish = finish;
    csv_file_dump fifo_csv_dumper_680;
    csv_file_dump cstatus_csv_dumper_680;
    df_fifo_monitor fifo_monitor_680;
    df_fifo_intf fifo_intf_681(clock,reset);
    assign fifo_intf_681.rd_en = AESL_inst_myproject.layer2_out_680_U.if_read & AESL_inst_myproject.layer2_out_680_U.if_empty_n;
    assign fifo_intf_681.wr_en = AESL_inst_myproject.layer2_out_680_U.if_write & AESL_inst_myproject.layer2_out_680_U.if_full_n;
    assign fifo_intf_681.fifo_rd_block = 0;
    assign fifo_intf_681.fifo_wr_block = 0;
    assign fifo_intf_681.finish = finish;
    csv_file_dump fifo_csv_dumper_681;
    csv_file_dump cstatus_csv_dumper_681;
    df_fifo_monitor fifo_monitor_681;
    df_fifo_intf fifo_intf_682(clock,reset);
    assign fifo_intf_682.rd_en = AESL_inst_myproject.layer2_out_681_U.if_read & AESL_inst_myproject.layer2_out_681_U.if_empty_n;
    assign fifo_intf_682.wr_en = AESL_inst_myproject.layer2_out_681_U.if_write & AESL_inst_myproject.layer2_out_681_U.if_full_n;
    assign fifo_intf_682.fifo_rd_block = 0;
    assign fifo_intf_682.fifo_wr_block = 0;
    assign fifo_intf_682.finish = finish;
    csv_file_dump fifo_csv_dumper_682;
    csv_file_dump cstatus_csv_dumper_682;
    df_fifo_monitor fifo_monitor_682;
    df_fifo_intf fifo_intf_683(clock,reset);
    assign fifo_intf_683.rd_en = AESL_inst_myproject.layer2_out_682_U.if_read & AESL_inst_myproject.layer2_out_682_U.if_empty_n;
    assign fifo_intf_683.wr_en = AESL_inst_myproject.layer2_out_682_U.if_write & AESL_inst_myproject.layer2_out_682_U.if_full_n;
    assign fifo_intf_683.fifo_rd_block = 0;
    assign fifo_intf_683.fifo_wr_block = 0;
    assign fifo_intf_683.finish = finish;
    csv_file_dump fifo_csv_dumper_683;
    csv_file_dump cstatus_csv_dumper_683;
    df_fifo_monitor fifo_monitor_683;
    df_fifo_intf fifo_intf_684(clock,reset);
    assign fifo_intf_684.rd_en = AESL_inst_myproject.layer2_out_683_U.if_read & AESL_inst_myproject.layer2_out_683_U.if_empty_n;
    assign fifo_intf_684.wr_en = AESL_inst_myproject.layer2_out_683_U.if_write & AESL_inst_myproject.layer2_out_683_U.if_full_n;
    assign fifo_intf_684.fifo_rd_block = 0;
    assign fifo_intf_684.fifo_wr_block = 0;
    assign fifo_intf_684.finish = finish;
    csv_file_dump fifo_csv_dumper_684;
    csv_file_dump cstatus_csv_dumper_684;
    df_fifo_monitor fifo_monitor_684;
    df_fifo_intf fifo_intf_685(clock,reset);
    assign fifo_intf_685.rd_en = AESL_inst_myproject.layer2_out_684_U.if_read & AESL_inst_myproject.layer2_out_684_U.if_empty_n;
    assign fifo_intf_685.wr_en = AESL_inst_myproject.layer2_out_684_U.if_write & AESL_inst_myproject.layer2_out_684_U.if_full_n;
    assign fifo_intf_685.fifo_rd_block = 0;
    assign fifo_intf_685.fifo_wr_block = 0;
    assign fifo_intf_685.finish = finish;
    csv_file_dump fifo_csv_dumper_685;
    csv_file_dump cstatus_csv_dumper_685;
    df_fifo_monitor fifo_monitor_685;
    df_fifo_intf fifo_intf_686(clock,reset);
    assign fifo_intf_686.rd_en = AESL_inst_myproject.layer2_out_685_U.if_read & AESL_inst_myproject.layer2_out_685_U.if_empty_n;
    assign fifo_intf_686.wr_en = AESL_inst_myproject.layer2_out_685_U.if_write & AESL_inst_myproject.layer2_out_685_U.if_full_n;
    assign fifo_intf_686.fifo_rd_block = 0;
    assign fifo_intf_686.fifo_wr_block = 0;
    assign fifo_intf_686.finish = finish;
    csv_file_dump fifo_csv_dumper_686;
    csv_file_dump cstatus_csv_dumper_686;
    df_fifo_monitor fifo_monitor_686;
    df_fifo_intf fifo_intf_687(clock,reset);
    assign fifo_intf_687.rd_en = AESL_inst_myproject.layer2_out_686_U.if_read & AESL_inst_myproject.layer2_out_686_U.if_empty_n;
    assign fifo_intf_687.wr_en = AESL_inst_myproject.layer2_out_686_U.if_write & AESL_inst_myproject.layer2_out_686_U.if_full_n;
    assign fifo_intf_687.fifo_rd_block = 0;
    assign fifo_intf_687.fifo_wr_block = 0;
    assign fifo_intf_687.finish = finish;
    csv_file_dump fifo_csv_dumper_687;
    csv_file_dump cstatus_csv_dumper_687;
    df_fifo_monitor fifo_monitor_687;
    df_fifo_intf fifo_intf_688(clock,reset);
    assign fifo_intf_688.rd_en = AESL_inst_myproject.layer2_out_687_U.if_read & AESL_inst_myproject.layer2_out_687_U.if_empty_n;
    assign fifo_intf_688.wr_en = AESL_inst_myproject.layer2_out_687_U.if_write & AESL_inst_myproject.layer2_out_687_U.if_full_n;
    assign fifo_intf_688.fifo_rd_block = 0;
    assign fifo_intf_688.fifo_wr_block = 0;
    assign fifo_intf_688.finish = finish;
    csv_file_dump fifo_csv_dumper_688;
    csv_file_dump cstatus_csv_dumper_688;
    df_fifo_monitor fifo_monitor_688;
    df_fifo_intf fifo_intf_689(clock,reset);
    assign fifo_intf_689.rd_en = AESL_inst_myproject.layer2_out_688_U.if_read & AESL_inst_myproject.layer2_out_688_U.if_empty_n;
    assign fifo_intf_689.wr_en = AESL_inst_myproject.layer2_out_688_U.if_write & AESL_inst_myproject.layer2_out_688_U.if_full_n;
    assign fifo_intf_689.fifo_rd_block = 0;
    assign fifo_intf_689.fifo_wr_block = 0;
    assign fifo_intf_689.finish = finish;
    csv_file_dump fifo_csv_dumper_689;
    csv_file_dump cstatus_csv_dumper_689;
    df_fifo_monitor fifo_monitor_689;
    df_fifo_intf fifo_intf_690(clock,reset);
    assign fifo_intf_690.rd_en = AESL_inst_myproject.layer2_out_689_U.if_read & AESL_inst_myproject.layer2_out_689_U.if_empty_n;
    assign fifo_intf_690.wr_en = AESL_inst_myproject.layer2_out_689_U.if_write & AESL_inst_myproject.layer2_out_689_U.if_full_n;
    assign fifo_intf_690.fifo_rd_block = 0;
    assign fifo_intf_690.fifo_wr_block = 0;
    assign fifo_intf_690.finish = finish;
    csv_file_dump fifo_csv_dumper_690;
    csv_file_dump cstatus_csv_dumper_690;
    df_fifo_monitor fifo_monitor_690;
    df_fifo_intf fifo_intf_691(clock,reset);
    assign fifo_intf_691.rd_en = AESL_inst_myproject.layer2_out_690_U.if_read & AESL_inst_myproject.layer2_out_690_U.if_empty_n;
    assign fifo_intf_691.wr_en = AESL_inst_myproject.layer2_out_690_U.if_write & AESL_inst_myproject.layer2_out_690_U.if_full_n;
    assign fifo_intf_691.fifo_rd_block = 0;
    assign fifo_intf_691.fifo_wr_block = 0;
    assign fifo_intf_691.finish = finish;
    csv_file_dump fifo_csv_dumper_691;
    csv_file_dump cstatus_csv_dumper_691;
    df_fifo_monitor fifo_monitor_691;
    df_fifo_intf fifo_intf_692(clock,reset);
    assign fifo_intf_692.rd_en = AESL_inst_myproject.layer2_out_691_U.if_read & AESL_inst_myproject.layer2_out_691_U.if_empty_n;
    assign fifo_intf_692.wr_en = AESL_inst_myproject.layer2_out_691_U.if_write & AESL_inst_myproject.layer2_out_691_U.if_full_n;
    assign fifo_intf_692.fifo_rd_block = 0;
    assign fifo_intf_692.fifo_wr_block = 0;
    assign fifo_intf_692.finish = finish;
    csv_file_dump fifo_csv_dumper_692;
    csv_file_dump cstatus_csv_dumper_692;
    df_fifo_monitor fifo_monitor_692;
    df_fifo_intf fifo_intf_693(clock,reset);
    assign fifo_intf_693.rd_en = AESL_inst_myproject.layer2_out_692_U.if_read & AESL_inst_myproject.layer2_out_692_U.if_empty_n;
    assign fifo_intf_693.wr_en = AESL_inst_myproject.layer2_out_692_U.if_write & AESL_inst_myproject.layer2_out_692_U.if_full_n;
    assign fifo_intf_693.fifo_rd_block = 0;
    assign fifo_intf_693.fifo_wr_block = 0;
    assign fifo_intf_693.finish = finish;
    csv_file_dump fifo_csv_dumper_693;
    csv_file_dump cstatus_csv_dumper_693;
    df_fifo_monitor fifo_monitor_693;
    df_fifo_intf fifo_intf_694(clock,reset);
    assign fifo_intf_694.rd_en = AESL_inst_myproject.layer2_out_693_U.if_read & AESL_inst_myproject.layer2_out_693_U.if_empty_n;
    assign fifo_intf_694.wr_en = AESL_inst_myproject.layer2_out_693_U.if_write & AESL_inst_myproject.layer2_out_693_U.if_full_n;
    assign fifo_intf_694.fifo_rd_block = 0;
    assign fifo_intf_694.fifo_wr_block = 0;
    assign fifo_intf_694.finish = finish;
    csv_file_dump fifo_csv_dumper_694;
    csv_file_dump cstatus_csv_dumper_694;
    df_fifo_monitor fifo_monitor_694;
    df_fifo_intf fifo_intf_695(clock,reset);
    assign fifo_intf_695.rd_en = AESL_inst_myproject.layer2_out_694_U.if_read & AESL_inst_myproject.layer2_out_694_U.if_empty_n;
    assign fifo_intf_695.wr_en = AESL_inst_myproject.layer2_out_694_U.if_write & AESL_inst_myproject.layer2_out_694_U.if_full_n;
    assign fifo_intf_695.fifo_rd_block = 0;
    assign fifo_intf_695.fifo_wr_block = 0;
    assign fifo_intf_695.finish = finish;
    csv_file_dump fifo_csv_dumper_695;
    csv_file_dump cstatus_csv_dumper_695;
    df_fifo_monitor fifo_monitor_695;
    df_fifo_intf fifo_intf_696(clock,reset);
    assign fifo_intf_696.rd_en = AESL_inst_myproject.layer2_out_695_U.if_read & AESL_inst_myproject.layer2_out_695_U.if_empty_n;
    assign fifo_intf_696.wr_en = AESL_inst_myproject.layer2_out_695_U.if_write & AESL_inst_myproject.layer2_out_695_U.if_full_n;
    assign fifo_intf_696.fifo_rd_block = 0;
    assign fifo_intf_696.fifo_wr_block = 0;
    assign fifo_intf_696.finish = finish;
    csv_file_dump fifo_csv_dumper_696;
    csv_file_dump cstatus_csv_dumper_696;
    df_fifo_monitor fifo_monitor_696;
    df_fifo_intf fifo_intf_697(clock,reset);
    assign fifo_intf_697.rd_en = AESL_inst_myproject.layer2_out_696_U.if_read & AESL_inst_myproject.layer2_out_696_U.if_empty_n;
    assign fifo_intf_697.wr_en = AESL_inst_myproject.layer2_out_696_U.if_write & AESL_inst_myproject.layer2_out_696_U.if_full_n;
    assign fifo_intf_697.fifo_rd_block = 0;
    assign fifo_intf_697.fifo_wr_block = 0;
    assign fifo_intf_697.finish = finish;
    csv_file_dump fifo_csv_dumper_697;
    csv_file_dump cstatus_csv_dumper_697;
    df_fifo_monitor fifo_monitor_697;
    df_fifo_intf fifo_intf_698(clock,reset);
    assign fifo_intf_698.rd_en = AESL_inst_myproject.layer2_out_697_U.if_read & AESL_inst_myproject.layer2_out_697_U.if_empty_n;
    assign fifo_intf_698.wr_en = AESL_inst_myproject.layer2_out_697_U.if_write & AESL_inst_myproject.layer2_out_697_U.if_full_n;
    assign fifo_intf_698.fifo_rd_block = 0;
    assign fifo_intf_698.fifo_wr_block = 0;
    assign fifo_intf_698.finish = finish;
    csv_file_dump fifo_csv_dumper_698;
    csv_file_dump cstatus_csv_dumper_698;
    df_fifo_monitor fifo_monitor_698;
    df_fifo_intf fifo_intf_699(clock,reset);
    assign fifo_intf_699.rd_en = AESL_inst_myproject.layer2_out_698_U.if_read & AESL_inst_myproject.layer2_out_698_U.if_empty_n;
    assign fifo_intf_699.wr_en = AESL_inst_myproject.layer2_out_698_U.if_write & AESL_inst_myproject.layer2_out_698_U.if_full_n;
    assign fifo_intf_699.fifo_rd_block = 0;
    assign fifo_intf_699.fifo_wr_block = 0;
    assign fifo_intf_699.finish = finish;
    csv_file_dump fifo_csv_dumper_699;
    csv_file_dump cstatus_csv_dumper_699;
    df_fifo_monitor fifo_monitor_699;
    df_fifo_intf fifo_intf_700(clock,reset);
    assign fifo_intf_700.rd_en = AESL_inst_myproject.layer2_out_699_U.if_read & AESL_inst_myproject.layer2_out_699_U.if_empty_n;
    assign fifo_intf_700.wr_en = AESL_inst_myproject.layer2_out_699_U.if_write & AESL_inst_myproject.layer2_out_699_U.if_full_n;
    assign fifo_intf_700.fifo_rd_block = 0;
    assign fifo_intf_700.fifo_wr_block = 0;
    assign fifo_intf_700.finish = finish;
    csv_file_dump fifo_csv_dumper_700;
    csv_file_dump cstatus_csv_dumper_700;
    df_fifo_monitor fifo_monitor_700;
    df_fifo_intf fifo_intf_701(clock,reset);
    assign fifo_intf_701.rd_en = AESL_inst_myproject.layer2_out_700_U.if_read & AESL_inst_myproject.layer2_out_700_U.if_empty_n;
    assign fifo_intf_701.wr_en = AESL_inst_myproject.layer2_out_700_U.if_write & AESL_inst_myproject.layer2_out_700_U.if_full_n;
    assign fifo_intf_701.fifo_rd_block = 0;
    assign fifo_intf_701.fifo_wr_block = 0;
    assign fifo_intf_701.finish = finish;
    csv_file_dump fifo_csv_dumper_701;
    csv_file_dump cstatus_csv_dumper_701;
    df_fifo_monitor fifo_monitor_701;
    df_fifo_intf fifo_intf_702(clock,reset);
    assign fifo_intf_702.rd_en = AESL_inst_myproject.layer2_out_701_U.if_read & AESL_inst_myproject.layer2_out_701_U.if_empty_n;
    assign fifo_intf_702.wr_en = AESL_inst_myproject.layer2_out_701_U.if_write & AESL_inst_myproject.layer2_out_701_U.if_full_n;
    assign fifo_intf_702.fifo_rd_block = 0;
    assign fifo_intf_702.fifo_wr_block = 0;
    assign fifo_intf_702.finish = finish;
    csv_file_dump fifo_csv_dumper_702;
    csv_file_dump cstatus_csv_dumper_702;
    df_fifo_monitor fifo_monitor_702;
    df_fifo_intf fifo_intf_703(clock,reset);
    assign fifo_intf_703.rd_en = AESL_inst_myproject.layer2_out_702_U.if_read & AESL_inst_myproject.layer2_out_702_U.if_empty_n;
    assign fifo_intf_703.wr_en = AESL_inst_myproject.layer2_out_702_U.if_write & AESL_inst_myproject.layer2_out_702_U.if_full_n;
    assign fifo_intf_703.fifo_rd_block = 0;
    assign fifo_intf_703.fifo_wr_block = 0;
    assign fifo_intf_703.finish = finish;
    csv_file_dump fifo_csv_dumper_703;
    csv_file_dump cstatus_csv_dumper_703;
    df_fifo_monitor fifo_monitor_703;
    df_fifo_intf fifo_intf_704(clock,reset);
    assign fifo_intf_704.rd_en = AESL_inst_myproject.layer2_out_703_U.if_read & AESL_inst_myproject.layer2_out_703_U.if_empty_n;
    assign fifo_intf_704.wr_en = AESL_inst_myproject.layer2_out_703_U.if_write & AESL_inst_myproject.layer2_out_703_U.if_full_n;
    assign fifo_intf_704.fifo_rd_block = 0;
    assign fifo_intf_704.fifo_wr_block = 0;
    assign fifo_intf_704.finish = finish;
    csv_file_dump fifo_csv_dumper_704;
    csv_file_dump cstatus_csv_dumper_704;
    df_fifo_monitor fifo_monitor_704;
    df_fifo_intf fifo_intf_705(clock,reset);
    assign fifo_intf_705.rd_en = AESL_inst_myproject.layer2_out_704_U.if_read & AESL_inst_myproject.layer2_out_704_U.if_empty_n;
    assign fifo_intf_705.wr_en = AESL_inst_myproject.layer2_out_704_U.if_write & AESL_inst_myproject.layer2_out_704_U.if_full_n;
    assign fifo_intf_705.fifo_rd_block = 0;
    assign fifo_intf_705.fifo_wr_block = 0;
    assign fifo_intf_705.finish = finish;
    csv_file_dump fifo_csv_dumper_705;
    csv_file_dump cstatus_csv_dumper_705;
    df_fifo_monitor fifo_monitor_705;
    df_fifo_intf fifo_intf_706(clock,reset);
    assign fifo_intf_706.rd_en = AESL_inst_myproject.layer2_out_705_U.if_read & AESL_inst_myproject.layer2_out_705_U.if_empty_n;
    assign fifo_intf_706.wr_en = AESL_inst_myproject.layer2_out_705_U.if_write & AESL_inst_myproject.layer2_out_705_U.if_full_n;
    assign fifo_intf_706.fifo_rd_block = 0;
    assign fifo_intf_706.fifo_wr_block = 0;
    assign fifo_intf_706.finish = finish;
    csv_file_dump fifo_csv_dumper_706;
    csv_file_dump cstatus_csv_dumper_706;
    df_fifo_monitor fifo_monitor_706;
    df_fifo_intf fifo_intf_707(clock,reset);
    assign fifo_intf_707.rd_en = AESL_inst_myproject.layer2_out_706_U.if_read & AESL_inst_myproject.layer2_out_706_U.if_empty_n;
    assign fifo_intf_707.wr_en = AESL_inst_myproject.layer2_out_706_U.if_write & AESL_inst_myproject.layer2_out_706_U.if_full_n;
    assign fifo_intf_707.fifo_rd_block = 0;
    assign fifo_intf_707.fifo_wr_block = 0;
    assign fifo_intf_707.finish = finish;
    csv_file_dump fifo_csv_dumper_707;
    csv_file_dump cstatus_csv_dumper_707;
    df_fifo_monitor fifo_monitor_707;
    df_fifo_intf fifo_intf_708(clock,reset);
    assign fifo_intf_708.rd_en = AESL_inst_myproject.layer2_out_707_U.if_read & AESL_inst_myproject.layer2_out_707_U.if_empty_n;
    assign fifo_intf_708.wr_en = AESL_inst_myproject.layer2_out_707_U.if_write & AESL_inst_myproject.layer2_out_707_U.if_full_n;
    assign fifo_intf_708.fifo_rd_block = 0;
    assign fifo_intf_708.fifo_wr_block = 0;
    assign fifo_intf_708.finish = finish;
    csv_file_dump fifo_csv_dumper_708;
    csv_file_dump cstatus_csv_dumper_708;
    df_fifo_monitor fifo_monitor_708;
    df_fifo_intf fifo_intf_709(clock,reset);
    assign fifo_intf_709.rd_en = AESL_inst_myproject.layer2_out_708_U.if_read & AESL_inst_myproject.layer2_out_708_U.if_empty_n;
    assign fifo_intf_709.wr_en = AESL_inst_myproject.layer2_out_708_U.if_write & AESL_inst_myproject.layer2_out_708_U.if_full_n;
    assign fifo_intf_709.fifo_rd_block = 0;
    assign fifo_intf_709.fifo_wr_block = 0;
    assign fifo_intf_709.finish = finish;
    csv_file_dump fifo_csv_dumper_709;
    csv_file_dump cstatus_csv_dumper_709;
    df_fifo_monitor fifo_monitor_709;
    df_fifo_intf fifo_intf_710(clock,reset);
    assign fifo_intf_710.rd_en = AESL_inst_myproject.layer2_out_709_U.if_read & AESL_inst_myproject.layer2_out_709_U.if_empty_n;
    assign fifo_intf_710.wr_en = AESL_inst_myproject.layer2_out_709_U.if_write & AESL_inst_myproject.layer2_out_709_U.if_full_n;
    assign fifo_intf_710.fifo_rd_block = 0;
    assign fifo_intf_710.fifo_wr_block = 0;
    assign fifo_intf_710.finish = finish;
    csv_file_dump fifo_csv_dumper_710;
    csv_file_dump cstatus_csv_dumper_710;
    df_fifo_monitor fifo_monitor_710;
    df_fifo_intf fifo_intf_711(clock,reset);
    assign fifo_intf_711.rd_en = AESL_inst_myproject.layer2_out_710_U.if_read & AESL_inst_myproject.layer2_out_710_U.if_empty_n;
    assign fifo_intf_711.wr_en = AESL_inst_myproject.layer2_out_710_U.if_write & AESL_inst_myproject.layer2_out_710_U.if_full_n;
    assign fifo_intf_711.fifo_rd_block = 0;
    assign fifo_intf_711.fifo_wr_block = 0;
    assign fifo_intf_711.finish = finish;
    csv_file_dump fifo_csv_dumper_711;
    csv_file_dump cstatus_csv_dumper_711;
    df_fifo_monitor fifo_monitor_711;
    df_fifo_intf fifo_intf_712(clock,reset);
    assign fifo_intf_712.rd_en = AESL_inst_myproject.layer2_out_711_U.if_read & AESL_inst_myproject.layer2_out_711_U.if_empty_n;
    assign fifo_intf_712.wr_en = AESL_inst_myproject.layer2_out_711_U.if_write & AESL_inst_myproject.layer2_out_711_U.if_full_n;
    assign fifo_intf_712.fifo_rd_block = 0;
    assign fifo_intf_712.fifo_wr_block = 0;
    assign fifo_intf_712.finish = finish;
    csv_file_dump fifo_csv_dumper_712;
    csv_file_dump cstatus_csv_dumper_712;
    df_fifo_monitor fifo_monitor_712;
    df_fifo_intf fifo_intf_713(clock,reset);
    assign fifo_intf_713.rd_en = AESL_inst_myproject.layer2_out_712_U.if_read & AESL_inst_myproject.layer2_out_712_U.if_empty_n;
    assign fifo_intf_713.wr_en = AESL_inst_myproject.layer2_out_712_U.if_write & AESL_inst_myproject.layer2_out_712_U.if_full_n;
    assign fifo_intf_713.fifo_rd_block = 0;
    assign fifo_intf_713.fifo_wr_block = 0;
    assign fifo_intf_713.finish = finish;
    csv_file_dump fifo_csv_dumper_713;
    csv_file_dump cstatus_csv_dumper_713;
    df_fifo_monitor fifo_monitor_713;
    df_fifo_intf fifo_intf_714(clock,reset);
    assign fifo_intf_714.rd_en = AESL_inst_myproject.layer2_out_713_U.if_read & AESL_inst_myproject.layer2_out_713_U.if_empty_n;
    assign fifo_intf_714.wr_en = AESL_inst_myproject.layer2_out_713_U.if_write & AESL_inst_myproject.layer2_out_713_U.if_full_n;
    assign fifo_intf_714.fifo_rd_block = 0;
    assign fifo_intf_714.fifo_wr_block = 0;
    assign fifo_intf_714.finish = finish;
    csv_file_dump fifo_csv_dumper_714;
    csv_file_dump cstatus_csv_dumper_714;
    df_fifo_monitor fifo_monitor_714;
    df_fifo_intf fifo_intf_715(clock,reset);
    assign fifo_intf_715.rd_en = AESL_inst_myproject.layer2_out_714_U.if_read & AESL_inst_myproject.layer2_out_714_U.if_empty_n;
    assign fifo_intf_715.wr_en = AESL_inst_myproject.layer2_out_714_U.if_write & AESL_inst_myproject.layer2_out_714_U.if_full_n;
    assign fifo_intf_715.fifo_rd_block = 0;
    assign fifo_intf_715.fifo_wr_block = 0;
    assign fifo_intf_715.finish = finish;
    csv_file_dump fifo_csv_dumper_715;
    csv_file_dump cstatus_csv_dumper_715;
    df_fifo_monitor fifo_monitor_715;
    df_fifo_intf fifo_intf_716(clock,reset);
    assign fifo_intf_716.rd_en = AESL_inst_myproject.layer2_out_715_U.if_read & AESL_inst_myproject.layer2_out_715_U.if_empty_n;
    assign fifo_intf_716.wr_en = AESL_inst_myproject.layer2_out_715_U.if_write & AESL_inst_myproject.layer2_out_715_U.if_full_n;
    assign fifo_intf_716.fifo_rd_block = 0;
    assign fifo_intf_716.fifo_wr_block = 0;
    assign fifo_intf_716.finish = finish;
    csv_file_dump fifo_csv_dumper_716;
    csv_file_dump cstatus_csv_dumper_716;
    df_fifo_monitor fifo_monitor_716;
    df_fifo_intf fifo_intf_717(clock,reset);
    assign fifo_intf_717.rd_en = AESL_inst_myproject.layer2_out_716_U.if_read & AESL_inst_myproject.layer2_out_716_U.if_empty_n;
    assign fifo_intf_717.wr_en = AESL_inst_myproject.layer2_out_716_U.if_write & AESL_inst_myproject.layer2_out_716_U.if_full_n;
    assign fifo_intf_717.fifo_rd_block = 0;
    assign fifo_intf_717.fifo_wr_block = 0;
    assign fifo_intf_717.finish = finish;
    csv_file_dump fifo_csv_dumper_717;
    csv_file_dump cstatus_csv_dumper_717;
    df_fifo_monitor fifo_monitor_717;
    df_fifo_intf fifo_intf_718(clock,reset);
    assign fifo_intf_718.rd_en = AESL_inst_myproject.layer2_out_717_U.if_read & AESL_inst_myproject.layer2_out_717_U.if_empty_n;
    assign fifo_intf_718.wr_en = AESL_inst_myproject.layer2_out_717_U.if_write & AESL_inst_myproject.layer2_out_717_U.if_full_n;
    assign fifo_intf_718.fifo_rd_block = 0;
    assign fifo_intf_718.fifo_wr_block = 0;
    assign fifo_intf_718.finish = finish;
    csv_file_dump fifo_csv_dumper_718;
    csv_file_dump cstatus_csv_dumper_718;
    df_fifo_monitor fifo_monitor_718;
    df_fifo_intf fifo_intf_719(clock,reset);
    assign fifo_intf_719.rd_en = AESL_inst_myproject.layer2_out_718_U.if_read & AESL_inst_myproject.layer2_out_718_U.if_empty_n;
    assign fifo_intf_719.wr_en = AESL_inst_myproject.layer2_out_718_U.if_write & AESL_inst_myproject.layer2_out_718_U.if_full_n;
    assign fifo_intf_719.fifo_rd_block = 0;
    assign fifo_intf_719.fifo_wr_block = 0;
    assign fifo_intf_719.finish = finish;
    csv_file_dump fifo_csv_dumper_719;
    csv_file_dump cstatus_csv_dumper_719;
    df_fifo_monitor fifo_monitor_719;
    df_fifo_intf fifo_intf_720(clock,reset);
    assign fifo_intf_720.rd_en = AESL_inst_myproject.layer2_out_719_U.if_read & AESL_inst_myproject.layer2_out_719_U.if_empty_n;
    assign fifo_intf_720.wr_en = AESL_inst_myproject.layer2_out_719_U.if_write & AESL_inst_myproject.layer2_out_719_U.if_full_n;
    assign fifo_intf_720.fifo_rd_block = 0;
    assign fifo_intf_720.fifo_wr_block = 0;
    assign fifo_intf_720.finish = finish;
    csv_file_dump fifo_csv_dumper_720;
    csv_file_dump cstatus_csv_dumper_720;
    df_fifo_monitor fifo_monitor_720;
    df_fifo_intf fifo_intf_721(clock,reset);
    assign fifo_intf_721.rd_en = AESL_inst_myproject.layer2_out_720_U.if_read & AESL_inst_myproject.layer2_out_720_U.if_empty_n;
    assign fifo_intf_721.wr_en = AESL_inst_myproject.layer2_out_720_U.if_write & AESL_inst_myproject.layer2_out_720_U.if_full_n;
    assign fifo_intf_721.fifo_rd_block = 0;
    assign fifo_intf_721.fifo_wr_block = 0;
    assign fifo_intf_721.finish = finish;
    csv_file_dump fifo_csv_dumper_721;
    csv_file_dump cstatus_csv_dumper_721;
    df_fifo_monitor fifo_monitor_721;
    df_fifo_intf fifo_intf_722(clock,reset);
    assign fifo_intf_722.rd_en = AESL_inst_myproject.layer2_out_721_U.if_read & AESL_inst_myproject.layer2_out_721_U.if_empty_n;
    assign fifo_intf_722.wr_en = AESL_inst_myproject.layer2_out_721_U.if_write & AESL_inst_myproject.layer2_out_721_U.if_full_n;
    assign fifo_intf_722.fifo_rd_block = 0;
    assign fifo_intf_722.fifo_wr_block = 0;
    assign fifo_intf_722.finish = finish;
    csv_file_dump fifo_csv_dumper_722;
    csv_file_dump cstatus_csv_dumper_722;
    df_fifo_monitor fifo_monitor_722;
    df_fifo_intf fifo_intf_723(clock,reset);
    assign fifo_intf_723.rd_en = AESL_inst_myproject.layer2_out_722_U.if_read & AESL_inst_myproject.layer2_out_722_U.if_empty_n;
    assign fifo_intf_723.wr_en = AESL_inst_myproject.layer2_out_722_U.if_write & AESL_inst_myproject.layer2_out_722_U.if_full_n;
    assign fifo_intf_723.fifo_rd_block = 0;
    assign fifo_intf_723.fifo_wr_block = 0;
    assign fifo_intf_723.finish = finish;
    csv_file_dump fifo_csv_dumper_723;
    csv_file_dump cstatus_csv_dumper_723;
    df_fifo_monitor fifo_monitor_723;
    df_fifo_intf fifo_intf_724(clock,reset);
    assign fifo_intf_724.rd_en = AESL_inst_myproject.layer2_out_723_U.if_read & AESL_inst_myproject.layer2_out_723_U.if_empty_n;
    assign fifo_intf_724.wr_en = AESL_inst_myproject.layer2_out_723_U.if_write & AESL_inst_myproject.layer2_out_723_U.if_full_n;
    assign fifo_intf_724.fifo_rd_block = 0;
    assign fifo_intf_724.fifo_wr_block = 0;
    assign fifo_intf_724.finish = finish;
    csv_file_dump fifo_csv_dumper_724;
    csv_file_dump cstatus_csv_dumper_724;
    df_fifo_monitor fifo_monitor_724;
    df_fifo_intf fifo_intf_725(clock,reset);
    assign fifo_intf_725.rd_en = AESL_inst_myproject.layer2_out_724_U.if_read & AESL_inst_myproject.layer2_out_724_U.if_empty_n;
    assign fifo_intf_725.wr_en = AESL_inst_myproject.layer2_out_724_U.if_write & AESL_inst_myproject.layer2_out_724_U.if_full_n;
    assign fifo_intf_725.fifo_rd_block = 0;
    assign fifo_intf_725.fifo_wr_block = 0;
    assign fifo_intf_725.finish = finish;
    csv_file_dump fifo_csv_dumper_725;
    csv_file_dump cstatus_csv_dumper_725;
    df_fifo_monitor fifo_monitor_725;
    df_fifo_intf fifo_intf_726(clock,reset);
    assign fifo_intf_726.rd_en = AESL_inst_myproject.layer2_out_725_U.if_read & AESL_inst_myproject.layer2_out_725_U.if_empty_n;
    assign fifo_intf_726.wr_en = AESL_inst_myproject.layer2_out_725_U.if_write & AESL_inst_myproject.layer2_out_725_U.if_full_n;
    assign fifo_intf_726.fifo_rd_block = 0;
    assign fifo_intf_726.fifo_wr_block = 0;
    assign fifo_intf_726.finish = finish;
    csv_file_dump fifo_csv_dumper_726;
    csv_file_dump cstatus_csv_dumper_726;
    df_fifo_monitor fifo_monitor_726;
    df_fifo_intf fifo_intf_727(clock,reset);
    assign fifo_intf_727.rd_en = AESL_inst_myproject.layer2_out_726_U.if_read & AESL_inst_myproject.layer2_out_726_U.if_empty_n;
    assign fifo_intf_727.wr_en = AESL_inst_myproject.layer2_out_726_U.if_write & AESL_inst_myproject.layer2_out_726_U.if_full_n;
    assign fifo_intf_727.fifo_rd_block = 0;
    assign fifo_intf_727.fifo_wr_block = 0;
    assign fifo_intf_727.finish = finish;
    csv_file_dump fifo_csv_dumper_727;
    csv_file_dump cstatus_csv_dumper_727;
    df_fifo_monitor fifo_monitor_727;
    df_fifo_intf fifo_intf_728(clock,reset);
    assign fifo_intf_728.rd_en = AESL_inst_myproject.layer2_out_727_U.if_read & AESL_inst_myproject.layer2_out_727_U.if_empty_n;
    assign fifo_intf_728.wr_en = AESL_inst_myproject.layer2_out_727_U.if_write & AESL_inst_myproject.layer2_out_727_U.if_full_n;
    assign fifo_intf_728.fifo_rd_block = 0;
    assign fifo_intf_728.fifo_wr_block = 0;
    assign fifo_intf_728.finish = finish;
    csv_file_dump fifo_csv_dumper_728;
    csv_file_dump cstatus_csv_dumper_728;
    df_fifo_monitor fifo_monitor_728;
    df_fifo_intf fifo_intf_729(clock,reset);
    assign fifo_intf_729.rd_en = AESL_inst_myproject.layer2_out_728_U.if_read & AESL_inst_myproject.layer2_out_728_U.if_empty_n;
    assign fifo_intf_729.wr_en = AESL_inst_myproject.layer2_out_728_U.if_write & AESL_inst_myproject.layer2_out_728_U.if_full_n;
    assign fifo_intf_729.fifo_rd_block = 0;
    assign fifo_intf_729.fifo_wr_block = 0;
    assign fifo_intf_729.finish = finish;
    csv_file_dump fifo_csv_dumper_729;
    csv_file_dump cstatus_csv_dumper_729;
    df_fifo_monitor fifo_monitor_729;
    df_fifo_intf fifo_intf_730(clock,reset);
    assign fifo_intf_730.rd_en = AESL_inst_myproject.layer2_out_729_U.if_read & AESL_inst_myproject.layer2_out_729_U.if_empty_n;
    assign fifo_intf_730.wr_en = AESL_inst_myproject.layer2_out_729_U.if_write & AESL_inst_myproject.layer2_out_729_U.if_full_n;
    assign fifo_intf_730.fifo_rd_block = 0;
    assign fifo_intf_730.fifo_wr_block = 0;
    assign fifo_intf_730.finish = finish;
    csv_file_dump fifo_csv_dumper_730;
    csv_file_dump cstatus_csv_dumper_730;
    df_fifo_monitor fifo_monitor_730;
    df_fifo_intf fifo_intf_731(clock,reset);
    assign fifo_intf_731.rd_en = AESL_inst_myproject.layer2_out_730_U.if_read & AESL_inst_myproject.layer2_out_730_U.if_empty_n;
    assign fifo_intf_731.wr_en = AESL_inst_myproject.layer2_out_730_U.if_write & AESL_inst_myproject.layer2_out_730_U.if_full_n;
    assign fifo_intf_731.fifo_rd_block = 0;
    assign fifo_intf_731.fifo_wr_block = 0;
    assign fifo_intf_731.finish = finish;
    csv_file_dump fifo_csv_dumper_731;
    csv_file_dump cstatus_csv_dumper_731;
    df_fifo_monitor fifo_monitor_731;
    df_fifo_intf fifo_intf_732(clock,reset);
    assign fifo_intf_732.rd_en = AESL_inst_myproject.layer2_out_731_U.if_read & AESL_inst_myproject.layer2_out_731_U.if_empty_n;
    assign fifo_intf_732.wr_en = AESL_inst_myproject.layer2_out_731_U.if_write & AESL_inst_myproject.layer2_out_731_U.if_full_n;
    assign fifo_intf_732.fifo_rd_block = 0;
    assign fifo_intf_732.fifo_wr_block = 0;
    assign fifo_intf_732.finish = finish;
    csv_file_dump fifo_csv_dumper_732;
    csv_file_dump cstatus_csv_dumper_732;
    df_fifo_monitor fifo_monitor_732;
    df_fifo_intf fifo_intf_733(clock,reset);
    assign fifo_intf_733.rd_en = AESL_inst_myproject.layer2_out_732_U.if_read & AESL_inst_myproject.layer2_out_732_U.if_empty_n;
    assign fifo_intf_733.wr_en = AESL_inst_myproject.layer2_out_732_U.if_write & AESL_inst_myproject.layer2_out_732_U.if_full_n;
    assign fifo_intf_733.fifo_rd_block = 0;
    assign fifo_intf_733.fifo_wr_block = 0;
    assign fifo_intf_733.finish = finish;
    csv_file_dump fifo_csv_dumper_733;
    csv_file_dump cstatus_csv_dumper_733;
    df_fifo_monitor fifo_monitor_733;
    df_fifo_intf fifo_intf_734(clock,reset);
    assign fifo_intf_734.rd_en = AESL_inst_myproject.layer2_out_733_U.if_read & AESL_inst_myproject.layer2_out_733_U.if_empty_n;
    assign fifo_intf_734.wr_en = AESL_inst_myproject.layer2_out_733_U.if_write & AESL_inst_myproject.layer2_out_733_U.if_full_n;
    assign fifo_intf_734.fifo_rd_block = 0;
    assign fifo_intf_734.fifo_wr_block = 0;
    assign fifo_intf_734.finish = finish;
    csv_file_dump fifo_csv_dumper_734;
    csv_file_dump cstatus_csv_dumper_734;
    df_fifo_monitor fifo_monitor_734;
    df_fifo_intf fifo_intf_735(clock,reset);
    assign fifo_intf_735.rd_en = AESL_inst_myproject.layer2_out_734_U.if_read & AESL_inst_myproject.layer2_out_734_U.if_empty_n;
    assign fifo_intf_735.wr_en = AESL_inst_myproject.layer2_out_734_U.if_write & AESL_inst_myproject.layer2_out_734_U.if_full_n;
    assign fifo_intf_735.fifo_rd_block = 0;
    assign fifo_intf_735.fifo_wr_block = 0;
    assign fifo_intf_735.finish = finish;
    csv_file_dump fifo_csv_dumper_735;
    csv_file_dump cstatus_csv_dumper_735;
    df_fifo_monitor fifo_monitor_735;
    df_fifo_intf fifo_intf_736(clock,reset);
    assign fifo_intf_736.rd_en = AESL_inst_myproject.layer2_out_735_U.if_read & AESL_inst_myproject.layer2_out_735_U.if_empty_n;
    assign fifo_intf_736.wr_en = AESL_inst_myproject.layer2_out_735_U.if_write & AESL_inst_myproject.layer2_out_735_U.if_full_n;
    assign fifo_intf_736.fifo_rd_block = 0;
    assign fifo_intf_736.fifo_wr_block = 0;
    assign fifo_intf_736.finish = finish;
    csv_file_dump fifo_csv_dumper_736;
    csv_file_dump cstatus_csv_dumper_736;
    df_fifo_monitor fifo_monitor_736;
    df_fifo_intf fifo_intf_737(clock,reset);
    assign fifo_intf_737.rd_en = AESL_inst_myproject.layer2_out_736_U.if_read & AESL_inst_myproject.layer2_out_736_U.if_empty_n;
    assign fifo_intf_737.wr_en = AESL_inst_myproject.layer2_out_736_U.if_write & AESL_inst_myproject.layer2_out_736_U.if_full_n;
    assign fifo_intf_737.fifo_rd_block = 0;
    assign fifo_intf_737.fifo_wr_block = 0;
    assign fifo_intf_737.finish = finish;
    csv_file_dump fifo_csv_dumper_737;
    csv_file_dump cstatus_csv_dumper_737;
    df_fifo_monitor fifo_monitor_737;
    df_fifo_intf fifo_intf_738(clock,reset);
    assign fifo_intf_738.rd_en = AESL_inst_myproject.layer2_out_737_U.if_read & AESL_inst_myproject.layer2_out_737_U.if_empty_n;
    assign fifo_intf_738.wr_en = AESL_inst_myproject.layer2_out_737_U.if_write & AESL_inst_myproject.layer2_out_737_U.if_full_n;
    assign fifo_intf_738.fifo_rd_block = 0;
    assign fifo_intf_738.fifo_wr_block = 0;
    assign fifo_intf_738.finish = finish;
    csv_file_dump fifo_csv_dumper_738;
    csv_file_dump cstatus_csv_dumper_738;
    df_fifo_monitor fifo_monitor_738;
    df_fifo_intf fifo_intf_739(clock,reset);
    assign fifo_intf_739.rd_en = AESL_inst_myproject.layer2_out_738_U.if_read & AESL_inst_myproject.layer2_out_738_U.if_empty_n;
    assign fifo_intf_739.wr_en = AESL_inst_myproject.layer2_out_738_U.if_write & AESL_inst_myproject.layer2_out_738_U.if_full_n;
    assign fifo_intf_739.fifo_rd_block = 0;
    assign fifo_intf_739.fifo_wr_block = 0;
    assign fifo_intf_739.finish = finish;
    csv_file_dump fifo_csv_dumper_739;
    csv_file_dump cstatus_csv_dumper_739;
    df_fifo_monitor fifo_monitor_739;
    df_fifo_intf fifo_intf_740(clock,reset);
    assign fifo_intf_740.rd_en = AESL_inst_myproject.layer2_out_739_U.if_read & AESL_inst_myproject.layer2_out_739_U.if_empty_n;
    assign fifo_intf_740.wr_en = AESL_inst_myproject.layer2_out_739_U.if_write & AESL_inst_myproject.layer2_out_739_U.if_full_n;
    assign fifo_intf_740.fifo_rd_block = 0;
    assign fifo_intf_740.fifo_wr_block = 0;
    assign fifo_intf_740.finish = finish;
    csv_file_dump fifo_csv_dumper_740;
    csv_file_dump cstatus_csv_dumper_740;
    df_fifo_monitor fifo_monitor_740;
    df_fifo_intf fifo_intf_741(clock,reset);
    assign fifo_intf_741.rd_en = AESL_inst_myproject.layer2_out_740_U.if_read & AESL_inst_myproject.layer2_out_740_U.if_empty_n;
    assign fifo_intf_741.wr_en = AESL_inst_myproject.layer2_out_740_U.if_write & AESL_inst_myproject.layer2_out_740_U.if_full_n;
    assign fifo_intf_741.fifo_rd_block = 0;
    assign fifo_intf_741.fifo_wr_block = 0;
    assign fifo_intf_741.finish = finish;
    csv_file_dump fifo_csv_dumper_741;
    csv_file_dump cstatus_csv_dumper_741;
    df_fifo_monitor fifo_monitor_741;
    df_fifo_intf fifo_intf_742(clock,reset);
    assign fifo_intf_742.rd_en = AESL_inst_myproject.layer2_out_741_U.if_read & AESL_inst_myproject.layer2_out_741_U.if_empty_n;
    assign fifo_intf_742.wr_en = AESL_inst_myproject.layer2_out_741_U.if_write & AESL_inst_myproject.layer2_out_741_U.if_full_n;
    assign fifo_intf_742.fifo_rd_block = 0;
    assign fifo_intf_742.fifo_wr_block = 0;
    assign fifo_intf_742.finish = finish;
    csv_file_dump fifo_csv_dumper_742;
    csv_file_dump cstatus_csv_dumper_742;
    df_fifo_monitor fifo_monitor_742;
    df_fifo_intf fifo_intf_743(clock,reset);
    assign fifo_intf_743.rd_en = AESL_inst_myproject.layer2_out_742_U.if_read & AESL_inst_myproject.layer2_out_742_U.if_empty_n;
    assign fifo_intf_743.wr_en = AESL_inst_myproject.layer2_out_742_U.if_write & AESL_inst_myproject.layer2_out_742_U.if_full_n;
    assign fifo_intf_743.fifo_rd_block = 0;
    assign fifo_intf_743.fifo_wr_block = 0;
    assign fifo_intf_743.finish = finish;
    csv_file_dump fifo_csv_dumper_743;
    csv_file_dump cstatus_csv_dumper_743;
    df_fifo_monitor fifo_monitor_743;
    df_fifo_intf fifo_intf_744(clock,reset);
    assign fifo_intf_744.rd_en = AESL_inst_myproject.layer2_out_743_U.if_read & AESL_inst_myproject.layer2_out_743_U.if_empty_n;
    assign fifo_intf_744.wr_en = AESL_inst_myproject.layer2_out_743_U.if_write & AESL_inst_myproject.layer2_out_743_U.if_full_n;
    assign fifo_intf_744.fifo_rd_block = 0;
    assign fifo_intf_744.fifo_wr_block = 0;
    assign fifo_intf_744.finish = finish;
    csv_file_dump fifo_csv_dumper_744;
    csv_file_dump cstatus_csv_dumper_744;
    df_fifo_monitor fifo_monitor_744;
    df_fifo_intf fifo_intf_745(clock,reset);
    assign fifo_intf_745.rd_en = AESL_inst_myproject.layer2_out_744_U.if_read & AESL_inst_myproject.layer2_out_744_U.if_empty_n;
    assign fifo_intf_745.wr_en = AESL_inst_myproject.layer2_out_744_U.if_write & AESL_inst_myproject.layer2_out_744_U.if_full_n;
    assign fifo_intf_745.fifo_rd_block = 0;
    assign fifo_intf_745.fifo_wr_block = 0;
    assign fifo_intf_745.finish = finish;
    csv_file_dump fifo_csv_dumper_745;
    csv_file_dump cstatus_csv_dumper_745;
    df_fifo_monitor fifo_monitor_745;
    df_fifo_intf fifo_intf_746(clock,reset);
    assign fifo_intf_746.rd_en = AESL_inst_myproject.layer2_out_745_U.if_read & AESL_inst_myproject.layer2_out_745_U.if_empty_n;
    assign fifo_intf_746.wr_en = AESL_inst_myproject.layer2_out_745_U.if_write & AESL_inst_myproject.layer2_out_745_U.if_full_n;
    assign fifo_intf_746.fifo_rd_block = 0;
    assign fifo_intf_746.fifo_wr_block = 0;
    assign fifo_intf_746.finish = finish;
    csv_file_dump fifo_csv_dumper_746;
    csv_file_dump cstatus_csv_dumper_746;
    df_fifo_monitor fifo_monitor_746;
    df_fifo_intf fifo_intf_747(clock,reset);
    assign fifo_intf_747.rd_en = AESL_inst_myproject.layer2_out_746_U.if_read & AESL_inst_myproject.layer2_out_746_U.if_empty_n;
    assign fifo_intf_747.wr_en = AESL_inst_myproject.layer2_out_746_U.if_write & AESL_inst_myproject.layer2_out_746_U.if_full_n;
    assign fifo_intf_747.fifo_rd_block = 0;
    assign fifo_intf_747.fifo_wr_block = 0;
    assign fifo_intf_747.finish = finish;
    csv_file_dump fifo_csv_dumper_747;
    csv_file_dump cstatus_csv_dumper_747;
    df_fifo_monitor fifo_monitor_747;
    df_fifo_intf fifo_intf_748(clock,reset);
    assign fifo_intf_748.rd_en = AESL_inst_myproject.layer2_out_747_U.if_read & AESL_inst_myproject.layer2_out_747_U.if_empty_n;
    assign fifo_intf_748.wr_en = AESL_inst_myproject.layer2_out_747_U.if_write & AESL_inst_myproject.layer2_out_747_U.if_full_n;
    assign fifo_intf_748.fifo_rd_block = 0;
    assign fifo_intf_748.fifo_wr_block = 0;
    assign fifo_intf_748.finish = finish;
    csv_file_dump fifo_csv_dumper_748;
    csv_file_dump cstatus_csv_dumper_748;
    df_fifo_monitor fifo_monitor_748;
    df_fifo_intf fifo_intf_749(clock,reset);
    assign fifo_intf_749.rd_en = AESL_inst_myproject.layer2_out_748_U.if_read & AESL_inst_myproject.layer2_out_748_U.if_empty_n;
    assign fifo_intf_749.wr_en = AESL_inst_myproject.layer2_out_748_U.if_write & AESL_inst_myproject.layer2_out_748_U.if_full_n;
    assign fifo_intf_749.fifo_rd_block = 0;
    assign fifo_intf_749.fifo_wr_block = 0;
    assign fifo_intf_749.finish = finish;
    csv_file_dump fifo_csv_dumper_749;
    csv_file_dump cstatus_csv_dumper_749;
    df_fifo_monitor fifo_monitor_749;
    df_fifo_intf fifo_intf_750(clock,reset);
    assign fifo_intf_750.rd_en = AESL_inst_myproject.layer2_out_749_U.if_read & AESL_inst_myproject.layer2_out_749_U.if_empty_n;
    assign fifo_intf_750.wr_en = AESL_inst_myproject.layer2_out_749_U.if_write & AESL_inst_myproject.layer2_out_749_U.if_full_n;
    assign fifo_intf_750.fifo_rd_block = 0;
    assign fifo_intf_750.fifo_wr_block = 0;
    assign fifo_intf_750.finish = finish;
    csv_file_dump fifo_csv_dumper_750;
    csv_file_dump cstatus_csv_dumper_750;
    df_fifo_monitor fifo_monitor_750;
    df_fifo_intf fifo_intf_751(clock,reset);
    assign fifo_intf_751.rd_en = AESL_inst_myproject.layer2_out_750_U.if_read & AESL_inst_myproject.layer2_out_750_U.if_empty_n;
    assign fifo_intf_751.wr_en = AESL_inst_myproject.layer2_out_750_U.if_write & AESL_inst_myproject.layer2_out_750_U.if_full_n;
    assign fifo_intf_751.fifo_rd_block = 0;
    assign fifo_intf_751.fifo_wr_block = 0;
    assign fifo_intf_751.finish = finish;
    csv_file_dump fifo_csv_dumper_751;
    csv_file_dump cstatus_csv_dumper_751;
    df_fifo_monitor fifo_monitor_751;
    df_fifo_intf fifo_intf_752(clock,reset);
    assign fifo_intf_752.rd_en = AESL_inst_myproject.layer2_out_751_U.if_read & AESL_inst_myproject.layer2_out_751_U.if_empty_n;
    assign fifo_intf_752.wr_en = AESL_inst_myproject.layer2_out_751_U.if_write & AESL_inst_myproject.layer2_out_751_U.if_full_n;
    assign fifo_intf_752.fifo_rd_block = 0;
    assign fifo_intf_752.fifo_wr_block = 0;
    assign fifo_intf_752.finish = finish;
    csv_file_dump fifo_csv_dumper_752;
    csv_file_dump cstatus_csv_dumper_752;
    df_fifo_monitor fifo_monitor_752;
    df_fifo_intf fifo_intf_753(clock,reset);
    assign fifo_intf_753.rd_en = AESL_inst_myproject.layer2_out_752_U.if_read & AESL_inst_myproject.layer2_out_752_U.if_empty_n;
    assign fifo_intf_753.wr_en = AESL_inst_myproject.layer2_out_752_U.if_write & AESL_inst_myproject.layer2_out_752_U.if_full_n;
    assign fifo_intf_753.fifo_rd_block = 0;
    assign fifo_intf_753.fifo_wr_block = 0;
    assign fifo_intf_753.finish = finish;
    csv_file_dump fifo_csv_dumper_753;
    csv_file_dump cstatus_csv_dumper_753;
    df_fifo_monitor fifo_monitor_753;
    df_fifo_intf fifo_intf_754(clock,reset);
    assign fifo_intf_754.rd_en = AESL_inst_myproject.layer2_out_753_U.if_read & AESL_inst_myproject.layer2_out_753_U.if_empty_n;
    assign fifo_intf_754.wr_en = AESL_inst_myproject.layer2_out_753_U.if_write & AESL_inst_myproject.layer2_out_753_U.if_full_n;
    assign fifo_intf_754.fifo_rd_block = 0;
    assign fifo_intf_754.fifo_wr_block = 0;
    assign fifo_intf_754.finish = finish;
    csv_file_dump fifo_csv_dumper_754;
    csv_file_dump cstatus_csv_dumper_754;
    df_fifo_monitor fifo_monitor_754;
    df_fifo_intf fifo_intf_755(clock,reset);
    assign fifo_intf_755.rd_en = AESL_inst_myproject.layer2_out_754_U.if_read & AESL_inst_myproject.layer2_out_754_U.if_empty_n;
    assign fifo_intf_755.wr_en = AESL_inst_myproject.layer2_out_754_U.if_write & AESL_inst_myproject.layer2_out_754_U.if_full_n;
    assign fifo_intf_755.fifo_rd_block = 0;
    assign fifo_intf_755.fifo_wr_block = 0;
    assign fifo_intf_755.finish = finish;
    csv_file_dump fifo_csv_dumper_755;
    csv_file_dump cstatus_csv_dumper_755;
    df_fifo_monitor fifo_monitor_755;
    df_fifo_intf fifo_intf_756(clock,reset);
    assign fifo_intf_756.rd_en = AESL_inst_myproject.layer2_out_755_U.if_read & AESL_inst_myproject.layer2_out_755_U.if_empty_n;
    assign fifo_intf_756.wr_en = AESL_inst_myproject.layer2_out_755_U.if_write & AESL_inst_myproject.layer2_out_755_U.if_full_n;
    assign fifo_intf_756.fifo_rd_block = 0;
    assign fifo_intf_756.fifo_wr_block = 0;
    assign fifo_intf_756.finish = finish;
    csv_file_dump fifo_csv_dumper_756;
    csv_file_dump cstatus_csv_dumper_756;
    df_fifo_monitor fifo_monitor_756;
    df_fifo_intf fifo_intf_757(clock,reset);
    assign fifo_intf_757.rd_en = AESL_inst_myproject.layer2_out_756_U.if_read & AESL_inst_myproject.layer2_out_756_U.if_empty_n;
    assign fifo_intf_757.wr_en = AESL_inst_myproject.layer2_out_756_U.if_write & AESL_inst_myproject.layer2_out_756_U.if_full_n;
    assign fifo_intf_757.fifo_rd_block = 0;
    assign fifo_intf_757.fifo_wr_block = 0;
    assign fifo_intf_757.finish = finish;
    csv_file_dump fifo_csv_dumper_757;
    csv_file_dump cstatus_csv_dumper_757;
    df_fifo_monitor fifo_monitor_757;
    df_fifo_intf fifo_intf_758(clock,reset);
    assign fifo_intf_758.rd_en = AESL_inst_myproject.layer2_out_757_U.if_read & AESL_inst_myproject.layer2_out_757_U.if_empty_n;
    assign fifo_intf_758.wr_en = AESL_inst_myproject.layer2_out_757_U.if_write & AESL_inst_myproject.layer2_out_757_U.if_full_n;
    assign fifo_intf_758.fifo_rd_block = 0;
    assign fifo_intf_758.fifo_wr_block = 0;
    assign fifo_intf_758.finish = finish;
    csv_file_dump fifo_csv_dumper_758;
    csv_file_dump cstatus_csv_dumper_758;
    df_fifo_monitor fifo_monitor_758;
    df_fifo_intf fifo_intf_759(clock,reset);
    assign fifo_intf_759.rd_en = AESL_inst_myproject.layer2_out_758_U.if_read & AESL_inst_myproject.layer2_out_758_U.if_empty_n;
    assign fifo_intf_759.wr_en = AESL_inst_myproject.layer2_out_758_U.if_write & AESL_inst_myproject.layer2_out_758_U.if_full_n;
    assign fifo_intf_759.fifo_rd_block = 0;
    assign fifo_intf_759.fifo_wr_block = 0;
    assign fifo_intf_759.finish = finish;
    csv_file_dump fifo_csv_dumper_759;
    csv_file_dump cstatus_csv_dumper_759;
    df_fifo_monitor fifo_monitor_759;
    df_fifo_intf fifo_intf_760(clock,reset);
    assign fifo_intf_760.rd_en = AESL_inst_myproject.layer2_out_759_U.if_read & AESL_inst_myproject.layer2_out_759_U.if_empty_n;
    assign fifo_intf_760.wr_en = AESL_inst_myproject.layer2_out_759_U.if_write & AESL_inst_myproject.layer2_out_759_U.if_full_n;
    assign fifo_intf_760.fifo_rd_block = 0;
    assign fifo_intf_760.fifo_wr_block = 0;
    assign fifo_intf_760.finish = finish;
    csv_file_dump fifo_csv_dumper_760;
    csv_file_dump cstatus_csv_dumper_760;
    df_fifo_monitor fifo_monitor_760;
    df_fifo_intf fifo_intf_761(clock,reset);
    assign fifo_intf_761.rd_en = AESL_inst_myproject.layer2_out_760_U.if_read & AESL_inst_myproject.layer2_out_760_U.if_empty_n;
    assign fifo_intf_761.wr_en = AESL_inst_myproject.layer2_out_760_U.if_write & AESL_inst_myproject.layer2_out_760_U.if_full_n;
    assign fifo_intf_761.fifo_rd_block = 0;
    assign fifo_intf_761.fifo_wr_block = 0;
    assign fifo_intf_761.finish = finish;
    csv_file_dump fifo_csv_dumper_761;
    csv_file_dump cstatus_csv_dumper_761;
    df_fifo_monitor fifo_monitor_761;
    df_fifo_intf fifo_intf_762(clock,reset);
    assign fifo_intf_762.rd_en = AESL_inst_myproject.layer2_out_761_U.if_read & AESL_inst_myproject.layer2_out_761_U.if_empty_n;
    assign fifo_intf_762.wr_en = AESL_inst_myproject.layer2_out_761_U.if_write & AESL_inst_myproject.layer2_out_761_U.if_full_n;
    assign fifo_intf_762.fifo_rd_block = 0;
    assign fifo_intf_762.fifo_wr_block = 0;
    assign fifo_intf_762.finish = finish;
    csv_file_dump fifo_csv_dumper_762;
    csv_file_dump cstatus_csv_dumper_762;
    df_fifo_monitor fifo_monitor_762;
    df_fifo_intf fifo_intf_763(clock,reset);
    assign fifo_intf_763.rd_en = AESL_inst_myproject.layer2_out_762_U.if_read & AESL_inst_myproject.layer2_out_762_U.if_empty_n;
    assign fifo_intf_763.wr_en = AESL_inst_myproject.layer2_out_762_U.if_write & AESL_inst_myproject.layer2_out_762_U.if_full_n;
    assign fifo_intf_763.fifo_rd_block = 0;
    assign fifo_intf_763.fifo_wr_block = 0;
    assign fifo_intf_763.finish = finish;
    csv_file_dump fifo_csv_dumper_763;
    csv_file_dump cstatus_csv_dumper_763;
    df_fifo_monitor fifo_monitor_763;
    df_fifo_intf fifo_intf_764(clock,reset);
    assign fifo_intf_764.rd_en = AESL_inst_myproject.layer2_out_763_U.if_read & AESL_inst_myproject.layer2_out_763_U.if_empty_n;
    assign fifo_intf_764.wr_en = AESL_inst_myproject.layer2_out_763_U.if_write & AESL_inst_myproject.layer2_out_763_U.if_full_n;
    assign fifo_intf_764.fifo_rd_block = 0;
    assign fifo_intf_764.fifo_wr_block = 0;
    assign fifo_intf_764.finish = finish;
    csv_file_dump fifo_csv_dumper_764;
    csv_file_dump cstatus_csv_dumper_764;
    df_fifo_monitor fifo_monitor_764;
    df_fifo_intf fifo_intf_765(clock,reset);
    assign fifo_intf_765.rd_en = AESL_inst_myproject.layer2_out_764_U.if_read & AESL_inst_myproject.layer2_out_764_U.if_empty_n;
    assign fifo_intf_765.wr_en = AESL_inst_myproject.layer2_out_764_U.if_write & AESL_inst_myproject.layer2_out_764_U.if_full_n;
    assign fifo_intf_765.fifo_rd_block = 0;
    assign fifo_intf_765.fifo_wr_block = 0;
    assign fifo_intf_765.finish = finish;
    csv_file_dump fifo_csv_dumper_765;
    csv_file_dump cstatus_csv_dumper_765;
    df_fifo_monitor fifo_monitor_765;
    df_fifo_intf fifo_intf_766(clock,reset);
    assign fifo_intf_766.rd_en = AESL_inst_myproject.layer2_out_765_U.if_read & AESL_inst_myproject.layer2_out_765_U.if_empty_n;
    assign fifo_intf_766.wr_en = AESL_inst_myproject.layer2_out_765_U.if_write & AESL_inst_myproject.layer2_out_765_U.if_full_n;
    assign fifo_intf_766.fifo_rd_block = 0;
    assign fifo_intf_766.fifo_wr_block = 0;
    assign fifo_intf_766.finish = finish;
    csv_file_dump fifo_csv_dumper_766;
    csv_file_dump cstatus_csv_dumper_766;
    df_fifo_monitor fifo_monitor_766;
    df_fifo_intf fifo_intf_767(clock,reset);
    assign fifo_intf_767.rd_en = AESL_inst_myproject.layer2_out_766_U.if_read & AESL_inst_myproject.layer2_out_766_U.if_empty_n;
    assign fifo_intf_767.wr_en = AESL_inst_myproject.layer2_out_766_U.if_write & AESL_inst_myproject.layer2_out_766_U.if_full_n;
    assign fifo_intf_767.fifo_rd_block = 0;
    assign fifo_intf_767.fifo_wr_block = 0;
    assign fifo_intf_767.finish = finish;
    csv_file_dump fifo_csv_dumper_767;
    csv_file_dump cstatus_csv_dumper_767;
    df_fifo_monitor fifo_monitor_767;
    df_fifo_intf fifo_intf_768(clock,reset);
    assign fifo_intf_768.rd_en = AESL_inst_myproject.layer2_out_767_U.if_read & AESL_inst_myproject.layer2_out_767_U.if_empty_n;
    assign fifo_intf_768.wr_en = AESL_inst_myproject.layer2_out_767_U.if_write & AESL_inst_myproject.layer2_out_767_U.if_full_n;
    assign fifo_intf_768.fifo_rd_block = 0;
    assign fifo_intf_768.fifo_wr_block = 0;
    assign fifo_intf_768.finish = finish;
    csv_file_dump fifo_csv_dumper_768;
    csv_file_dump cstatus_csv_dumper_768;
    df_fifo_monitor fifo_monitor_768;
    df_fifo_intf fifo_intf_769(clock,reset);
    assign fifo_intf_769.rd_en = AESL_inst_myproject.layer2_out_768_U.if_read & AESL_inst_myproject.layer2_out_768_U.if_empty_n;
    assign fifo_intf_769.wr_en = AESL_inst_myproject.layer2_out_768_U.if_write & AESL_inst_myproject.layer2_out_768_U.if_full_n;
    assign fifo_intf_769.fifo_rd_block = 0;
    assign fifo_intf_769.fifo_wr_block = 0;
    assign fifo_intf_769.finish = finish;
    csv_file_dump fifo_csv_dumper_769;
    csv_file_dump cstatus_csv_dumper_769;
    df_fifo_monitor fifo_monitor_769;
    df_fifo_intf fifo_intf_770(clock,reset);
    assign fifo_intf_770.rd_en = AESL_inst_myproject.layer2_out_769_U.if_read & AESL_inst_myproject.layer2_out_769_U.if_empty_n;
    assign fifo_intf_770.wr_en = AESL_inst_myproject.layer2_out_769_U.if_write & AESL_inst_myproject.layer2_out_769_U.if_full_n;
    assign fifo_intf_770.fifo_rd_block = 0;
    assign fifo_intf_770.fifo_wr_block = 0;
    assign fifo_intf_770.finish = finish;
    csv_file_dump fifo_csv_dumper_770;
    csv_file_dump cstatus_csv_dumper_770;
    df_fifo_monitor fifo_monitor_770;
    df_fifo_intf fifo_intf_771(clock,reset);
    assign fifo_intf_771.rd_en = AESL_inst_myproject.layer2_out_770_U.if_read & AESL_inst_myproject.layer2_out_770_U.if_empty_n;
    assign fifo_intf_771.wr_en = AESL_inst_myproject.layer2_out_770_U.if_write & AESL_inst_myproject.layer2_out_770_U.if_full_n;
    assign fifo_intf_771.fifo_rd_block = 0;
    assign fifo_intf_771.fifo_wr_block = 0;
    assign fifo_intf_771.finish = finish;
    csv_file_dump fifo_csv_dumper_771;
    csv_file_dump cstatus_csv_dumper_771;
    df_fifo_monitor fifo_monitor_771;
    df_fifo_intf fifo_intf_772(clock,reset);
    assign fifo_intf_772.rd_en = AESL_inst_myproject.layer2_out_771_U.if_read & AESL_inst_myproject.layer2_out_771_U.if_empty_n;
    assign fifo_intf_772.wr_en = AESL_inst_myproject.layer2_out_771_U.if_write & AESL_inst_myproject.layer2_out_771_U.if_full_n;
    assign fifo_intf_772.fifo_rd_block = 0;
    assign fifo_intf_772.fifo_wr_block = 0;
    assign fifo_intf_772.finish = finish;
    csv_file_dump fifo_csv_dumper_772;
    csv_file_dump cstatus_csv_dumper_772;
    df_fifo_monitor fifo_monitor_772;
    df_fifo_intf fifo_intf_773(clock,reset);
    assign fifo_intf_773.rd_en = AESL_inst_myproject.layer2_out_772_U.if_read & AESL_inst_myproject.layer2_out_772_U.if_empty_n;
    assign fifo_intf_773.wr_en = AESL_inst_myproject.layer2_out_772_U.if_write & AESL_inst_myproject.layer2_out_772_U.if_full_n;
    assign fifo_intf_773.fifo_rd_block = 0;
    assign fifo_intf_773.fifo_wr_block = 0;
    assign fifo_intf_773.finish = finish;
    csv_file_dump fifo_csv_dumper_773;
    csv_file_dump cstatus_csv_dumper_773;
    df_fifo_monitor fifo_monitor_773;
    df_fifo_intf fifo_intf_774(clock,reset);
    assign fifo_intf_774.rd_en = AESL_inst_myproject.layer2_out_773_U.if_read & AESL_inst_myproject.layer2_out_773_U.if_empty_n;
    assign fifo_intf_774.wr_en = AESL_inst_myproject.layer2_out_773_U.if_write & AESL_inst_myproject.layer2_out_773_U.if_full_n;
    assign fifo_intf_774.fifo_rd_block = 0;
    assign fifo_intf_774.fifo_wr_block = 0;
    assign fifo_intf_774.finish = finish;
    csv_file_dump fifo_csv_dumper_774;
    csv_file_dump cstatus_csv_dumper_774;
    df_fifo_monitor fifo_monitor_774;
    df_fifo_intf fifo_intf_775(clock,reset);
    assign fifo_intf_775.rd_en = AESL_inst_myproject.layer2_out_774_U.if_read & AESL_inst_myproject.layer2_out_774_U.if_empty_n;
    assign fifo_intf_775.wr_en = AESL_inst_myproject.layer2_out_774_U.if_write & AESL_inst_myproject.layer2_out_774_U.if_full_n;
    assign fifo_intf_775.fifo_rd_block = 0;
    assign fifo_intf_775.fifo_wr_block = 0;
    assign fifo_intf_775.finish = finish;
    csv_file_dump fifo_csv_dumper_775;
    csv_file_dump cstatus_csv_dumper_775;
    df_fifo_monitor fifo_monitor_775;
    df_fifo_intf fifo_intf_776(clock,reset);
    assign fifo_intf_776.rd_en = AESL_inst_myproject.layer2_out_775_U.if_read & AESL_inst_myproject.layer2_out_775_U.if_empty_n;
    assign fifo_intf_776.wr_en = AESL_inst_myproject.layer2_out_775_U.if_write & AESL_inst_myproject.layer2_out_775_U.if_full_n;
    assign fifo_intf_776.fifo_rd_block = 0;
    assign fifo_intf_776.fifo_wr_block = 0;
    assign fifo_intf_776.finish = finish;
    csv_file_dump fifo_csv_dumper_776;
    csv_file_dump cstatus_csv_dumper_776;
    df_fifo_monitor fifo_monitor_776;
    df_fifo_intf fifo_intf_777(clock,reset);
    assign fifo_intf_777.rd_en = AESL_inst_myproject.layer2_out_776_U.if_read & AESL_inst_myproject.layer2_out_776_U.if_empty_n;
    assign fifo_intf_777.wr_en = AESL_inst_myproject.layer2_out_776_U.if_write & AESL_inst_myproject.layer2_out_776_U.if_full_n;
    assign fifo_intf_777.fifo_rd_block = 0;
    assign fifo_intf_777.fifo_wr_block = 0;
    assign fifo_intf_777.finish = finish;
    csv_file_dump fifo_csv_dumper_777;
    csv_file_dump cstatus_csv_dumper_777;
    df_fifo_monitor fifo_monitor_777;
    df_fifo_intf fifo_intf_778(clock,reset);
    assign fifo_intf_778.rd_en = AESL_inst_myproject.layer2_out_777_U.if_read & AESL_inst_myproject.layer2_out_777_U.if_empty_n;
    assign fifo_intf_778.wr_en = AESL_inst_myproject.layer2_out_777_U.if_write & AESL_inst_myproject.layer2_out_777_U.if_full_n;
    assign fifo_intf_778.fifo_rd_block = 0;
    assign fifo_intf_778.fifo_wr_block = 0;
    assign fifo_intf_778.finish = finish;
    csv_file_dump fifo_csv_dumper_778;
    csv_file_dump cstatus_csv_dumper_778;
    df_fifo_monitor fifo_monitor_778;
    df_fifo_intf fifo_intf_779(clock,reset);
    assign fifo_intf_779.rd_en = AESL_inst_myproject.layer2_out_778_U.if_read & AESL_inst_myproject.layer2_out_778_U.if_empty_n;
    assign fifo_intf_779.wr_en = AESL_inst_myproject.layer2_out_778_U.if_write & AESL_inst_myproject.layer2_out_778_U.if_full_n;
    assign fifo_intf_779.fifo_rd_block = 0;
    assign fifo_intf_779.fifo_wr_block = 0;
    assign fifo_intf_779.finish = finish;
    csv_file_dump fifo_csv_dumper_779;
    csv_file_dump cstatus_csv_dumper_779;
    df_fifo_monitor fifo_monitor_779;
    df_fifo_intf fifo_intf_780(clock,reset);
    assign fifo_intf_780.rd_en = AESL_inst_myproject.layer2_out_779_U.if_read & AESL_inst_myproject.layer2_out_779_U.if_empty_n;
    assign fifo_intf_780.wr_en = AESL_inst_myproject.layer2_out_779_U.if_write & AESL_inst_myproject.layer2_out_779_U.if_full_n;
    assign fifo_intf_780.fifo_rd_block = 0;
    assign fifo_intf_780.fifo_wr_block = 0;
    assign fifo_intf_780.finish = finish;
    csv_file_dump fifo_csv_dumper_780;
    csv_file_dump cstatus_csv_dumper_780;
    df_fifo_monitor fifo_monitor_780;
    df_fifo_intf fifo_intf_781(clock,reset);
    assign fifo_intf_781.rd_en = AESL_inst_myproject.layer2_out_780_U.if_read & AESL_inst_myproject.layer2_out_780_U.if_empty_n;
    assign fifo_intf_781.wr_en = AESL_inst_myproject.layer2_out_780_U.if_write & AESL_inst_myproject.layer2_out_780_U.if_full_n;
    assign fifo_intf_781.fifo_rd_block = 0;
    assign fifo_intf_781.fifo_wr_block = 0;
    assign fifo_intf_781.finish = finish;
    csv_file_dump fifo_csv_dumper_781;
    csv_file_dump cstatus_csv_dumper_781;
    df_fifo_monitor fifo_monitor_781;
    df_fifo_intf fifo_intf_782(clock,reset);
    assign fifo_intf_782.rd_en = AESL_inst_myproject.layer2_out_781_U.if_read & AESL_inst_myproject.layer2_out_781_U.if_empty_n;
    assign fifo_intf_782.wr_en = AESL_inst_myproject.layer2_out_781_U.if_write & AESL_inst_myproject.layer2_out_781_U.if_full_n;
    assign fifo_intf_782.fifo_rd_block = 0;
    assign fifo_intf_782.fifo_wr_block = 0;
    assign fifo_intf_782.finish = finish;
    csv_file_dump fifo_csv_dumper_782;
    csv_file_dump cstatus_csv_dumper_782;
    df_fifo_monitor fifo_monitor_782;
    df_fifo_intf fifo_intf_783(clock,reset);
    assign fifo_intf_783.rd_en = AESL_inst_myproject.layer2_out_782_U.if_read & AESL_inst_myproject.layer2_out_782_U.if_empty_n;
    assign fifo_intf_783.wr_en = AESL_inst_myproject.layer2_out_782_U.if_write & AESL_inst_myproject.layer2_out_782_U.if_full_n;
    assign fifo_intf_783.fifo_rd_block = 0;
    assign fifo_intf_783.fifo_wr_block = 0;
    assign fifo_intf_783.finish = finish;
    csv_file_dump fifo_csv_dumper_783;
    csv_file_dump cstatus_csv_dumper_783;
    df_fifo_monitor fifo_monitor_783;
    df_fifo_intf fifo_intf_784(clock,reset);
    assign fifo_intf_784.rd_en = AESL_inst_myproject.layer2_out_783_U.if_read & AESL_inst_myproject.layer2_out_783_U.if_empty_n;
    assign fifo_intf_784.wr_en = AESL_inst_myproject.layer2_out_783_U.if_write & AESL_inst_myproject.layer2_out_783_U.if_full_n;
    assign fifo_intf_784.fifo_rd_block = 0;
    assign fifo_intf_784.fifo_wr_block = 0;
    assign fifo_intf_784.finish = finish;
    csv_file_dump fifo_csv_dumper_784;
    csv_file_dump cstatus_csv_dumper_784;
    df_fifo_monitor fifo_monitor_784;
    df_fifo_intf fifo_intf_785(clock,reset);
    assign fifo_intf_785.rd_en = AESL_inst_myproject.layer2_out_784_U.if_read & AESL_inst_myproject.layer2_out_784_U.if_empty_n;
    assign fifo_intf_785.wr_en = AESL_inst_myproject.layer2_out_784_U.if_write & AESL_inst_myproject.layer2_out_784_U.if_full_n;
    assign fifo_intf_785.fifo_rd_block = 0;
    assign fifo_intf_785.fifo_wr_block = 0;
    assign fifo_intf_785.finish = finish;
    csv_file_dump fifo_csv_dumper_785;
    csv_file_dump cstatus_csv_dumper_785;
    df_fifo_monitor fifo_monitor_785;
    df_fifo_intf fifo_intf_786(clock,reset);
    assign fifo_intf_786.rd_en = AESL_inst_myproject.layer2_out_785_U.if_read & AESL_inst_myproject.layer2_out_785_U.if_empty_n;
    assign fifo_intf_786.wr_en = AESL_inst_myproject.layer2_out_785_U.if_write & AESL_inst_myproject.layer2_out_785_U.if_full_n;
    assign fifo_intf_786.fifo_rd_block = 0;
    assign fifo_intf_786.fifo_wr_block = 0;
    assign fifo_intf_786.finish = finish;
    csv_file_dump fifo_csv_dumper_786;
    csv_file_dump cstatus_csv_dumper_786;
    df_fifo_monitor fifo_monitor_786;
    df_fifo_intf fifo_intf_787(clock,reset);
    assign fifo_intf_787.rd_en = AESL_inst_myproject.layer2_out_786_U.if_read & AESL_inst_myproject.layer2_out_786_U.if_empty_n;
    assign fifo_intf_787.wr_en = AESL_inst_myproject.layer2_out_786_U.if_write & AESL_inst_myproject.layer2_out_786_U.if_full_n;
    assign fifo_intf_787.fifo_rd_block = 0;
    assign fifo_intf_787.fifo_wr_block = 0;
    assign fifo_intf_787.finish = finish;
    csv_file_dump fifo_csv_dumper_787;
    csv_file_dump cstatus_csv_dumper_787;
    df_fifo_monitor fifo_monitor_787;
    df_fifo_intf fifo_intf_788(clock,reset);
    assign fifo_intf_788.rd_en = AESL_inst_myproject.layer2_out_787_U.if_read & AESL_inst_myproject.layer2_out_787_U.if_empty_n;
    assign fifo_intf_788.wr_en = AESL_inst_myproject.layer2_out_787_U.if_write & AESL_inst_myproject.layer2_out_787_U.if_full_n;
    assign fifo_intf_788.fifo_rd_block = 0;
    assign fifo_intf_788.fifo_wr_block = 0;
    assign fifo_intf_788.finish = finish;
    csv_file_dump fifo_csv_dumper_788;
    csv_file_dump cstatus_csv_dumper_788;
    df_fifo_monitor fifo_monitor_788;
    df_fifo_intf fifo_intf_789(clock,reset);
    assign fifo_intf_789.rd_en = AESL_inst_myproject.layer2_out_788_U.if_read & AESL_inst_myproject.layer2_out_788_U.if_empty_n;
    assign fifo_intf_789.wr_en = AESL_inst_myproject.layer2_out_788_U.if_write & AESL_inst_myproject.layer2_out_788_U.if_full_n;
    assign fifo_intf_789.fifo_rd_block = 0;
    assign fifo_intf_789.fifo_wr_block = 0;
    assign fifo_intf_789.finish = finish;
    csv_file_dump fifo_csv_dumper_789;
    csv_file_dump cstatus_csv_dumper_789;
    df_fifo_monitor fifo_monitor_789;
    df_fifo_intf fifo_intf_790(clock,reset);
    assign fifo_intf_790.rd_en = AESL_inst_myproject.layer2_out_789_U.if_read & AESL_inst_myproject.layer2_out_789_U.if_empty_n;
    assign fifo_intf_790.wr_en = AESL_inst_myproject.layer2_out_789_U.if_write & AESL_inst_myproject.layer2_out_789_U.if_full_n;
    assign fifo_intf_790.fifo_rd_block = 0;
    assign fifo_intf_790.fifo_wr_block = 0;
    assign fifo_intf_790.finish = finish;
    csv_file_dump fifo_csv_dumper_790;
    csv_file_dump cstatus_csv_dumper_790;
    df_fifo_monitor fifo_monitor_790;
    df_fifo_intf fifo_intf_791(clock,reset);
    assign fifo_intf_791.rd_en = AESL_inst_myproject.layer2_out_790_U.if_read & AESL_inst_myproject.layer2_out_790_U.if_empty_n;
    assign fifo_intf_791.wr_en = AESL_inst_myproject.layer2_out_790_U.if_write & AESL_inst_myproject.layer2_out_790_U.if_full_n;
    assign fifo_intf_791.fifo_rd_block = 0;
    assign fifo_intf_791.fifo_wr_block = 0;
    assign fifo_intf_791.finish = finish;
    csv_file_dump fifo_csv_dumper_791;
    csv_file_dump cstatus_csv_dumper_791;
    df_fifo_monitor fifo_monitor_791;
    df_fifo_intf fifo_intf_792(clock,reset);
    assign fifo_intf_792.rd_en = AESL_inst_myproject.layer2_out_791_U.if_read & AESL_inst_myproject.layer2_out_791_U.if_empty_n;
    assign fifo_intf_792.wr_en = AESL_inst_myproject.layer2_out_791_U.if_write & AESL_inst_myproject.layer2_out_791_U.if_full_n;
    assign fifo_intf_792.fifo_rd_block = 0;
    assign fifo_intf_792.fifo_wr_block = 0;
    assign fifo_intf_792.finish = finish;
    csv_file_dump fifo_csv_dumper_792;
    csv_file_dump cstatus_csv_dumper_792;
    df_fifo_monitor fifo_monitor_792;
    df_fifo_intf fifo_intf_793(clock,reset);
    assign fifo_intf_793.rd_en = AESL_inst_myproject.layer2_out_792_U.if_read & AESL_inst_myproject.layer2_out_792_U.if_empty_n;
    assign fifo_intf_793.wr_en = AESL_inst_myproject.layer2_out_792_U.if_write & AESL_inst_myproject.layer2_out_792_U.if_full_n;
    assign fifo_intf_793.fifo_rd_block = 0;
    assign fifo_intf_793.fifo_wr_block = 0;
    assign fifo_intf_793.finish = finish;
    csv_file_dump fifo_csv_dumper_793;
    csv_file_dump cstatus_csv_dumper_793;
    df_fifo_monitor fifo_monitor_793;
    df_fifo_intf fifo_intf_794(clock,reset);
    assign fifo_intf_794.rd_en = AESL_inst_myproject.layer2_out_793_U.if_read & AESL_inst_myproject.layer2_out_793_U.if_empty_n;
    assign fifo_intf_794.wr_en = AESL_inst_myproject.layer2_out_793_U.if_write & AESL_inst_myproject.layer2_out_793_U.if_full_n;
    assign fifo_intf_794.fifo_rd_block = 0;
    assign fifo_intf_794.fifo_wr_block = 0;
    assign fifo_intf_794.finish = finish;
    csv_file_dump fifo_csv_dumper_794;
    csv_file_dump cstatus_csv_dumper_794;
    df_fifo_monitor fifo_monitor_794;
    df_fifo_intf fifo_intf_795(clock,reset);
    assign fifo_intf_795.rd_en = AESL_inst_myproject.layer2_out_794_U.if_read & AESL_inst_myproject.layer2_out_794_U.if_empty_n;
    assign fifo_intf_795.wr_en = AESL_inst_myproject.layer2_out_794_U.if_write & AESL_inst_myproject.layer2_out_794_U.if_full_n;
    assign fifo_intf_795.fifo_rd_block = 0;
    assign fifo_intf_795.fifo_wr_block = 0;
    assign fifo_intf_795.finish = finish;
    csv_file_dump fifo_csv_dumper_795;
    csv_file_dump cstatus_csv_dumper_795;
    df_fifo_monitor fifo_monitor_795;
    df_fifo_intf fifo_intf_796(clock,reset);
    assign fifo_intf_796.rd_en = AESL_inst_myproject.layer2_out_795_U.if_read & AESL_inst_myproject.layer2_out_795_U.if_empty_n;
    assign fifo_intf_796.wr_en = AESL_inst_myproject.layer2_out_795_U.if_write & AESL_inst_myproject.layer2_out_795_U.if_full_n;
    assign fifo_intf_796.fifo_rd_block = 0;
    assign fifo_intf_796.fifo_wr_block = 0;
    assign fifo_intf_796.finish = finish;
    csv_file_dump fifo_csv_dumper_796;
    csv_file_dump cstatus_csv_dumper_796;
    df_fifo_monitor fifo_monitor_796;
    df_fifo_intf fifo_intf_797(clock,reset);
    assign fifo_intf_797.rd_en = AESL_inst_myproject.layer2_out_796_U.if_read & AESL_inst_myproject.layer2_out_796_U.if_empty_n;
    assign fifo_intf_797.wr_en = AESL_inst_myproject.layer2_out_796_U.if_write & AESL_inst_myproject.layer2_out_796_U.if_full_n;
    assign fifo_intf_797.fifo_rd_block = 0;
    assign fifo_intf_797.fifo_wr_block = 0;
    assign fifo_intf_797.finish = finish;
    csv_file_dump fifo_csv_dumper_797;
    csv_file_dump cstatus_csv_dumper_797;
    df_fifo_monitor fifo_monitor_797;
    df_fifo_intf fifo_intf_798(clock,reset);
    assign fifo_intf_798.rd_en = AESL_inst_myproject.layer2_out_797_U.if_read & AESL_inst_myproject.layer2_out_797_U.if_empty_n;
    assign fifo_intf_798.wr_en = AESL_inst_myproject.layer2_out_797_U.if_write & AESL_inst_myproject.layer2_out_797_U.if_full_n;
    assign fifo_intf_798.fifo_rd_block = 0;
    assign fifo_intf_798.fifo_wr_block = 0;
    assign fifo_intf_798.finish = finish;
    csv_file_dump fifo_csv_dumper_798;
    csv_file_dump cstatus_csv_dumper_798;
    df_fifo_monitor fifo_monitor_798;
    df_fifo_intf fifo_intf_799(clock,reset);
    assign fifo_intf_799.rd_en = AESL_inst_myproject.layer2_out_798_U.if_read & AESL_inst_myproject.layer2_out_798_U.if_empty_n;
    assign fifo_intf_799.wr_en = AESL_inst_myproject.layer2_out_798_U.if_write & AESL_inst_myproject.layer2_out_798_U.if_full_n;
    assign fifo_intf_799.fifo_rd_block = 0;
    assign fifo_intf_799.fifo_wr_block = 0;
    assign fifo_intf_799.finish = finish;
    csv_file_dump fifo_csv_dumper_799;
    csv_file_dump cstatus_csv_dumper_799;
    df_fifo_monitor fifo_monitor_799;
    df_fifo_intf fifo_intf_800(clock,reset);
    assign fifo_intf_800.rd_en = AESL_inst_myproject.layer2_out_799_U.if_read & AESL_inst_myproject.layer2_out_799_U.if_empty_n;
    assign fifo_intf_800.wr_en = AESL_inst_myproject.layer2_out_799_U.if_write & AESL_inst_myproject.layer2_out_799_U.if_full_n;
    assign fifo_intf_800.fifo_rd_block = 0;
    assign fifo_intf_800.fifo_wr_block = 0;
    assign fifo_intf_800.finish = finish;
    csv_file_dump fifo_csv_dumper_800;
    csv_file_dump cstatus_csv_dumper_800;
    df_fifo_monitor fifo_monitor_800;
    df_fifo_intf fifo_intf_801(clock,reset);
    assign fifo_intf_801.rd_en = AESL_inst_myproject.layer2_out_800_U.if_read & AESL_inst_myproject.layer2_out_800_U.if_empty_n;
    assign fifo_intf_801.wr_en = AESL_inst_myproject.layer2_out_800_U.if_write & AESL_inst_myproject.layer2_out_800_U.if_full_n;
    assign fifo_intf_801.fifo_rd_block = 0;
    assign fifo_intf_801.fifo_wr_block = 0;
    assign fifo_intf_801.finish = finish;
    csv_file_dump fifo_csv_dumper_801;
    csv_file_dump cstatus_csv_dumper_801;
    df_fifo_monitor fifo_monitor_801;
    df_fifo_intf fifo_intf_802(clock,reset);
    assign fifo_intf_802.rd_en = AESL_inst_myproject.layer2_out_801_U.if_read & AESL_inst_myproject.layer2_out_801_U.if_empty_n;
    assign fifo_intf_802.wr_en = AESL_inst_myproject.layer2_out_801_U.if_write & AESL_inst_myproject.layer2_out_801_U.if_full_n;
    assign fifo_intf_802.fifo_rd_block = 0;
    assign fifo_intf_802.fifo_wr_block = 0;
    assign fifo_intf_802.finish = finish;
    csv_file_dump fifo_csv_dumper_802;
    csv_file_dump cstatus_csv_dumper_802;
    df_fifo_monitor fifo_monitor_802;
    df_fifo_intf fifo_intf_803(clock,reset);
    assign fifo_intf_803.rd_en = AESL_inst_myproject.layer2_out_802_U.if_read & AESL_inst_myproject.layer2_out_802_U.if_empty_n;
    assign fifo_intf_803.wr_en = AESL_inst_myproject.layer2_out_802_U.if_write & AESL_inst_myproject.layer2_out_802_U.if_full_n;
    assign fifo_intf_803.fifo_rd_block = 0;
    assign fifo_intf_803.fifo_wr_block = 0;
    assign fifo_intf_803.finish = finish;
    csv_file_dump fifo_csv_dumper_803;
    csv_file_dump cstatus_csv_dumper_803;
    df_fifo_monitor fifo_monitor_803;
    df_fifo_intf fifo_intf_804(clock,reset);
    assign fifo_intf_804.rd_en = AESL_inst_myproject.layer2_out_803_U.if_read & AESL_inst_myproject.layer2_out_803_U.if_empty_n;
    assign fifo_intf_804.wr_en = AESL_inst_myproject.layer2_out_803_U.if_write & AESL_inst_myproject.layer2_out_803_U.if_full_n;
    assign fifo_intf_804.fifo_rd_block = 0;
    assign fifo_intf_804.fifo_wr_block = 0;
    assign fifo_intf_804.finish = finish;
    csv_file_dump fifo_csv_dumper_804;
    csv_file_dump cstatus_csv_dumper_804;
    df_fifo_monitor fifo_monitor_804;
    df_fifo_intf fifo_intf_805(clock,reset);
    assign fifo_intf_805.rd_en = AESL_inst_myproject.layer2_out_804_U.if_read & AESL_inst_myproject.layer2_out_804_U.if_empty_n;
    assign fifo_intf_805.wr_en = AESL_inst_myproject.layer2_out_804_U.if_write & AESL_inst_myproject.layer2_out_804_U.if_full_n;
    assign fifo_intf_805.fifo_rd_block = 0;
    assign fifo_intf_805.fifo_wr_block = 0;
    assign fifo_intf_805.finish = finish;
    csv_file_dump fifo_csv_dumper_805;
    csv_file_dump cstatus_csv_dumper_805;
    df_fifo_monitor fifo_monitor_805;
    df_fifo_intf fifo_intf_806(clock,reset);
    assign fifo_intf_806.rd_en = AESL_inst_myproject.layer2_out_805_U.if_read & AESL_inst_myproject.layer2_out_805_U.if_empty_n;
    assign fifo_intf_806.wr_en = AESL_inst_myproject.layer2_out_805_U.if_write & AESL_inst_myproject.layer2_out_805_U.if_full_n;
    assign fifo_intf_806.fifo_rd_block = 0;
    assign fifo_intf_806.fifo_wr_block = 0;
    assign fifo_intf_806.finish = finish;
    csv_file_dump fifo_csv_dumper_806;
    csv_file_dump cstatus_csv_dumper_806;
    df_fifo_monitor fifo_monitor_806;
    df_fifo_intf fifo_intf_807(clock,reset);
    assign fifo_intf_807.rd_en = AESL_inst_myproject.layer2_out_806_U.if_read & AESL_inst_myproject.layer2_out_806_U.if_empty_n;
    assign fifo_intf_807.wr_en = AESL_inst_myproject.layer2_out_806_U.if_write & AESL_inst_myproject.layer2_out_806_U.if_full_n;
    assign fifo_intf_807.fifo_rd_block = 0;
    assign fifo_intf_807.fifo_wr_block = 0;
    assign fifo_intf_807.finish = finish;
    csv_file_dump fifo_csv_dumper_807;
    csv_file_dump cstatus_csv_dumper_807;
    df_fifo_monitor fifo_monitor_807;
    df_fifo_intf fifo_intf_808(clock,reset);
    assign fifo_intf_808.rd_en = AESL_inst_myproject.layer2_out_807_U.if_read & AESL_inst_myproject.layer2_out_807_U.if_empty_n;
    assign fifo_intf_808.wr_en = AESL_inst_myproject.layer2_out_807_U.if_write & AESL_inst_myproject.layer2_out_807_U.if_full_n;
    assign fifo_intf_808.fifo_rd_block = 0;
    assign fifo_intf_808.fifo_wr_block = 0;
    assign fifo_intf_808.finish = finish;
    csv_file_dump fifo_csv_dumper_808;
    csv_file_dump cstatus_csv_dumper_808;
    df_fifo_monitor fifo_monitor_808;
    df_fifo_intf fifo_intf_809(clock,reset);
    assign fifo_intf_809.rd_en = AESL_inst_myproject.layer2_out_808_U.if_read & AESL_inst_myproject.layer2_out_808_U.if_empty_n;
    assign fifo_intf_809.wr_en = AESL_inst_myproject.layer2_out_808_U.if_write & AESL_inst_myproject.layer2_out_808_U.if_full_n;
    assign fifo_intf_809.fifo_rd_block = 0;
    assign fifo_intf_809.fifo_wr_block = 0;
    assign fifo_intf_809.finish = finish;
    csv_file_dump fifo_csv_dumper_809;
    csv_file_dump cstatus_csv_dumper_809;
    df_fifo_monitor fifo_monitor_809;
    df_fifo_intf fifo_intf_810(clock,reset);
    assign fifo_intf_810.rd_en = AESL_inst_myproject.layer2_out_809_U.if_read & AESL_inst_myproject.layer2_out_809_U.if_empty_n;
    assign fifo_intf_810.wr_en = AESL_inst_myproject.layer2_out_809_U.if_write & AESL_inst_myproject.layer2_out_809_U.if_full_n;
    assign fifo_intf_810.fifo_rd_block = 0;
    assign fifo_intf_810.fifo_wr_block = 0;
    assign fifo_intf_810.finish = finish;
    csv_file_dump fifo_csv_dumper_810;
    csv_file_dump cstatus_csv_dumper_810;
    df_fifo_monitor fifo_monitor_810;
    df_fifo_intf fifo_intf_811(clock,reset);
    assign fifo_intf_811.rd_en = AESL_inst_myproject.layer2_out_810_U.if_read & AESL_inst_myproject.layer2_out_810_U.if_empty_n;
    assign fifo_intf_811.wr_en = AESL_inst_myproject.layer2_out_810_U.if_write & AESL_inst_myproject.layer2_out_810_U.if_full_n;
    assign fifo_intf_811.fifo_rd_block = 0;
    assign fifo_intf_811.fifo_wr_block = 0;
    assign fifo_intf_811.finish = finish;
    csv_file_dump fifo_csv_dumper_811;
    csv_file_dump cstatus_csv_dumper_811;
    df_fifo_monitor fifo_monitor_811;
    df_fifo_intf fifo_intf_812(clock,reset);
    assign fifo_intf_812.rd_en = AESL_inst_myproject.layer2_out_811_U.if_read & AESL_inst_myproject.layer2_out_811_U.if_empty_n;
    assign fifo_intf_812.wr_en = AESL_inst_myproject.layer2_out_811_U.if_write & AESL_inst_myproject.layer2_out_811_U.if_full_n;
    assign fifo_intf_812.fifo_rd_block = 0;
    assign fifo_intf_812.fifo_wr_block = 0;
    assign fifo_intf_812.finish = finish;
    csv_file_dump fifo_csv_dumper_812;
    csv_file_dump cstatus_csv_dumper_812;
    df_fifo_monitor fifo_monitor_812;
    df_fifo_intf fifo_intf_813(clock,reset);
    assign fifo_intf_813.rd_en = AESL_inst_myproject.layer2_out_812_U.if_read & AESL_inst_myproject.layer2_out_812_U.if_empty_n;
    assign fifo_intf_813.wr_en = AESL_inst_myproject.layer2_out_812_U.if_write & AESL_inst_myproject.layer2_out_812_U.if_full_n;
    assign fifo_intf_813.fifo_rd_block = 0;
    assign fifo_intf_813.fifo_wr_block = 0;
    assign fifo_intf_813.finish = finish;
    csv_file_dump fifo_csv_dumper_813;
    csv_file_dump cstatus_csv_dumper_813;
    df_fifo_monitor fifo_monitor_813;
    df_fifo_intf fifo_intf_814(clock,reset);
    assign fifo_intf_814.rd_en = AESL_inst_myproject.layer2_out_813_U.if_read & AESL_inst_myproject.layer2_out_813_U.if_empty_n;
    assign fifo_intf_814.wr_en = AESL_inst_myproject.layer2_out_813_U.if_write & AESL_inst_myproject.layer2_out_813_U.if_full_n;
    assign fifo_intf_814.fifo_rd_block = 0;
    assign fifo_intf_814.fifo_wr_block = 0;
    assign fifo_intf_814.finish = finish;
    csv_file_dump fifo_csv_dumper_814;
    csv_file_dump cstatus_csv_dumper_814;
    df_fifo_monitor fifo_monitor_814;
    df_fifo_intf fifo_intf_815(clock,reset);
    assign fifo_intf_815.rd_en = AESL_inst_myproject.layer2_out_814_U.if_read & AESL_inst_myproject.layer2_out_814_U.if_empty_n;
    assign fifo_intf_815.wr_en = AESL_inst_myproject.layer2_out_814_U.if_write & AESL_inst_myproject.layer2_out_814_U.if_full_n;
    assign fifo_intf_815.fifo_rd_block = 0;
    assign fifo_intf_815.fifo_wr_block = 0;
    assign fifo_intf_815.finish = finish;
    csv_file_dump fifo_csv_dumper_815;
    csv_file_dump cstatus_csv_dumper_815;
    df_fifo_monitor fifo_monitor_815;
    df_fifo_intf fifo_intf_816(clock,reset);
    assign fifo_intf_816.rd_en = AESL_inst_myproject.layer2_out_815_U.if_read & AESL_inst_myproject.layer2_out_815_U.if_empty_n;
    assign fifo_intf_816.wr_en = AESL_inst_myproject.layer2_out_815_U.if_write & AESL_inst_myproject.layer2_out_815_U.if_full_n;
    assign fifo_intf_816.fifo_rd_block = 0;
    assign fifo_intf_816.fifo_wr_block = 0;
    assign fifo_intf_816.finish = finish;
    csv_file_dump fifo_csv_dumper_816;
    csv_file_dump cstatus_csv_dumper_816;
    df_fifo_monitor fifo_monitor_816;
    df_fifo_intf fifo_intf_817(clock,reset);
    assign fifo_intf_817.rd_en = AESL_inst_myproject.layer2_out_816_U.if_read & AESL_inst_myproject.layer2_out_816_U.if_empty_n;
    assign fifo_intf_817.wr_en = AESL_inst_myproject.layer2_out_816_U.if_write & AESL_inst_myproject.layer2_out_816_U.if_full_n;
    assign fifo_intf_817.fifo_rd_block = 0;
    assign fifo_intf_817.fifo_wr_block = 0;
    assign fifo_intf_817.finish = finish;
    csv_file_dump fifo_csv_dumper_817;
    csv_file_dump cstatus_csv_dumper_817;
    df_fifo_monitor fifo_monitor_817;
    df_fifo_intf fifo_intf_818(clock,reset);
    assign fifo_intf_818.rd_en = AESL_inst_myproject.layer2_out_817_U.if_read & AESL_inst_myproject.layer2_out_817_U.if_empty_n;
    assign fifo_intf_818.wr_en = AESL_inst_myproject.layer2_out_817_U.if_write & AESL_inst_myproject.layer2_out_817_U.if_full_n;
    assign fifo_intf_818.fifo_rd_block = 0;
    assign fifo_intf_818.fifo_wr_block = 0;
    assign fifo_intf_818.finish = finish;
    csv_file_dump fifo_csv_dumper_818;
    csv_file_dump cstatus_csv_dumper_818;
    df_fifo_monitor fifo_monitor_818;
    df_fifo_intf fifo_intf_819(clock,reset);
    assign fifo_intf_819.rd_en = AESL_inst_myproject.layer2_out_818_U.if_read & AESL_inst_myproject.layer2_out_818_U.if_empty_n;
    assign fifo_intf_819.wr_en = AESL_inst_myproject.layer2_out_818_U.if_write & AESL_inst_myproject.layer2_out_818_U.if_full_n;
    assign fifo_intf_819.fifo_rd_block = 0;
    assign fifo_intf_819.fifo_wr_block = 0;
    assign fifo_intf_819.finish = finish;
    csv_file_dump fifo_csv_dumper_819;
    csv_file_dump cstatus_csv_dumper_819;
    df_fifo_monitor fifo_monitor_819;
    df_fifo_intf fifo_intf_820(clock,reset);
    assign fifo_intf_820.rd_en = AESL_inst_myproject.layer2_out_819_U.if_read & AESL_inst_myproject.layer2_out_819_U.if_empty_n;
    assign fifo_intf_820.wr_en = AESL_inst_myproject.layer2_out_819_U.if_write & AESL_inst_myproject.layer2_out_819_U.if_full_n;
    assign fifo_intf_820.fifo_rd_block = 0;
    assign fifo_intf_820.fifo_wr_block = 0;
    assign fifo_intf_820.finish = finish;
    csv_file_dump fifo_csv_dumper_820;
    csv_file_dump cstatus_csv_dumper_820;
    df_fifo_monitor fifo_monitor_820;
    df_fifo_intf fifo_intf_821(clock,reset);
    assign fifo_intf_821.rd_en = AESL_inst_myproject.layer2_out_820_U.if_read & AESL_inst_myproject.layer2_out_820_U.if_empty_n;
    assign fifo_intf_821.wr_en = AESL_inst_myproject.layer2_out_820_U.if_write & AESL_inst_myproject.layer2_out_820_U.if_full_n;
    assign fifo_intf_821.fifo_rd_block = 0;
    assign fifo_intf_821.fifo_wr_block = 0;
    assign fifo_intf_821.finish = finish;
    csv_file_dump fifo_csv_dumper_821;
    csv_file_dump cstatus_csv_dumper_821;
    df_fifo_monitor fifo_monitor_821;
    df_fifo_intf fifo_intf_822(clock,reset);
    assign fifo_intf_822.rd_en = AESL_inst_myproject.layer2_out_821_U.if_read & AESL_inst_myproject.layer2_out_821_U.if_empty_n;
    assign fifo_intf_822.wr_en = AESL_inst_myproject.layer2_out_821_U.if_write & AESL_inst_myproject.layer2_out_821_U.if_full_n;
    assign fifo_intf_822.fifo_rd_block = 0;
    assign fifo_intf_822.fifo_wr_block = 0;
    assign fifo_intf_822.finish = finish;
    csv_file_dump fifo_csv_dumper_822;
    csv_file_dump cstatus_csv_dumper_822;
    df_fifo_monitor fifo_monitor_822;
    df_fifo_intf fifo_intf_823(clock,reset);
    assign fifo_intf_823.rd_en = AESL_inst_myproject.layer2_out_822_U.if_read & AESL_inst_myproject.layer2_out_822_U.if_empty_n;
    assign fifo_intf_823.wr_en = AESL_inst_myproject.layer2_out_822_U.if_write & AESL_inst_myproject.layer2_out_822_U.if_full_n;
    assign fifo_intf_823.fifo_rd_block = 0;
    assign fifo_intf_823.fifo_wr_block = 0;
    assign fifo_intf_823.finish = finish;
    csv_file_dump fifo_csv_dumper_823;
    csv_file_dump cstatus_csv_dumper_823;
    df_fifo_monitor fifo_monitor_823;
    df_fifo_intf fifo_intf_824(clock,reset);
    assign fifo_intf_824.rd_en = AESL_inst_myproject.layer2_out_823_U.if_read & AESL_inst_myproject.layer2_out_823_U.if_empty_n;
    assign fifo_intf_824.wr_en = AESL_inst_myproject.layer2_out_823_U.if_write & AESL_inst_myproject.layer2_out_823_U.if_full_n;
    assign fifo_intf_824.fifo_rd_block = 0;
    assign fifo_intf_824.fifo_wr_block = 0;
    assign fifo_intf_824.finish = finish;
    csv_file_dump fifo_csv_dumper_824;
    csv_file_dump cstatus_csv_dumper_824;
    df_fifo_monitor fifo_monitor_824;
    df_fifo_intf fifo_intf_825(clock,reset);
    assign fifo_intf_825.rd_en = AESL_inst_myproject.layer2_out_824_U.if_read & AESL_inst_myproject.layer2_out_824_U.if_empty_n;
    assign fifo_intf_825.wr_en = AESL_inst_myproject.layer2_out_824_U.if_write & AESL_inst_myproject.layer2_out_824_U.if_full_n;
    assign fifo_intf_825.fifo_rd_block = 0;
    assign fifo_intf_825.fifo_wr_block = 0;
    assign fifo_intf_825.finish = finish;
    csv_file_dump fifo_csv_dumper_825;
    csv_file_dump cstatus_csv_dumper_825;
    df_fifo_monitor fifo_monitor_825;
    df_fifo_intf fifo_intf_826(clock,reset);
    assign fifo_intf_826.rd_en = AESL_inst_myproject.layer2_out_825_U.if_read & AESL_inst_myproject.layer2_out_825_U.if_empty_n;
    assign fifo_intf_826.wr_en = AESL_inst_myproject.layer2_out_825_U.if_write & AESL_inst_myproject.layer2_out_825_U.if_full_n;
    assign fifo_intf_826.fifo_rd_block = 0;
    assign fifo_intf_826.fifo_wr_block = 0;
    assign fifo_intf_826.finish = finish;
    csv_file_dump fifo_csv_dumper_826;
    csv_file_dump cstatus_csv_dumper_826;
    df_fifo_monitor fifo_monitor_826;
    df_fifo_intf fifo_intf_827(clock,reset);
    assign fifo_intf_827.rd_en = AESL_inst_myproject.layer2_out_826_U.if_read & AESL_inst_myproject.layer2_out_826_U.if_empty_n;
    assign fifo_intf_827.wr_en = AESL_inst_myproject.layer2_out_826_U.if_write & AESL_inst_myproject.layer2_out_826_U.if_full_n;
    assign fifo_intf_827.fifo_rd_block = 0;
    assign fifo_intf_827.fifo_wr_block = 0;
    assign fifo_intf_827.finish = finish;
    csv_file_dump fifo_csv_dumper_827;
    csv_file_dump cstatus_csv_dumper_827;
    df_fifo_monitor fifo_monitor_827;
    df_fifo_intf fifo_intf_828(clock,reset);
    assign fifo_intf_828.rd_en = AESL_inst_myproject.layer2_out_827_U.if_read & AESL_inst_myproject.layer2_out_827_U.if_empty_n;
    assign fifo_intf_828.wr_en = AESL_inst_myproject.layer2_out_827_U.if_write & AESL_inst_myproject.layer2_out_827_U.if_full_n;
    assign fifo_intf_828.fifo_rd_block = 0;
    assign fifo_intf_828.fifo_wr_block = 0;
    assign fifo_intf_828.finish = finish;
    csv_file_dump fifo_csv_dumper_828;
    csv_file_dump cstatus_csv_dumper_828;
    df_fifo_monitor fifo_monitor_828;
    df_fifo_intf fifo_intf_829(clock,reset);
    assign fifo_intf_829.rd_en = AESL_inst_myproject.layer2_out_828_U.if_read & AESL_inst_myproject.layer2_out_828_U.if_empty_n;
    assign fifo_intf_829.wr_en = AESL_inst_myproject.layer2_out_828_U.if_write & AESL_inst_myproject.layer2_out_828_U.if_full_n;
    assign fifo_intf_829.fifo_rd_block = 0;
    assign fifo_intf_829.fifo_wr_block = 0;
    assign fifo_intf_829.finish = finish;
    csv_file_dump fifo_csv_dumper_829;
    csv_file_dump cstatus_csv_dumper_829;
    df_fifo_monitor fifo_monitor_829;
    df_fifo_intf fifo_intf_830(clock,reset);
    assign fifo_intf_830.rd_en = AESL_inst_myproject.layer2_out_829_U.if_read & AESL_inst_myproject.layer2_out_829_U.if_empty_n;
    assign fifo_intf_830.wr_en = AESL_inst_myproject.layer2_out_829_U.if_write & AESL_inst_myproject.layer2_out_829_U.if_full_n;
    assign fifo_intf_830.fifo_rd_block = 0;
    assign fifo_intf_830.fifo_wr_block = 0;
    assign fifo_intf_830.finish = finish;
    csv_file_dump fifo_csv_dumper_830;
    csv_file_dump cstatus_csv_dumper_830;
    df_fifo_monitor fifo_monitor_830;
    df_fifo_intf fifo_intf_831(clock,reset);
    assign fifo_intf_831.rd_en = AESL_inst_myproject.layer2_out_830_U.if_read & AESL_inst_myproject.layer2_out_830_U.if_empty_n;
    assign fifo_intf_831.wr_en = AESL_inst_myproject.layer2_out_830_U.if_write & AESL_inst_myproject.layer2_out_830_U.if_full_n;
    assign fifo_intf_831.fifo_rd_block = 0;
    assign fifo_intf_831.fifo_wr_block = 0;
    assign fifo_intf_831.finish = finish;
    csv_file_dump fifo_csv_dumper_831;
    csv_file_dump cstatus_csv_dumper_831;
    df_fifo_monitor fifo_monitor_831;
    df_fifo_intf fifo_intf_832(clock,reset);
    assign fifo_intf_832.rd_en = AESL_inst_myproject.layer2_out_831_U.if_read & AESL_inst_myproject.layer2_out_831_U.if_empty_n;
    assign fifo_intf_832.wr_en = AESL_inst_myproject.layer2_out_831_U.if_write & AESL_inst_myproject.layer2_out_831_U.if_full_n;
    assign fifo_intf_832.fifo_rd_block = 0;
    assign fifo_intf_832.fifo_wr_block = 0;
    assign fifo_intf_832.finish = finish;
    csv_file_dump fifo_csv_dumper_832;
    csv_file_dump cstatus_csv_dumper_832;
    df_fifo_monitor fifo_monitor_832;
    df_fifo_intf fifo_intf_833(clock,reset);
    assign fifo_intf_833.rd_en = AESL_inst_myproject.layer2_out_832_U.if_read & AESL_inst_myproject.layer2_out_832_U.if_empty_n;
    assign fifo_intf_833.wr_en = AESL_inst_myproject.layer2_out_832_U.if_write & AESL_inst_myproject.layer2_out_832_U.if_full_n;
    assign fifo_intf_833.fifo_rd_block = 0;
    assign fifo_intf_833.fifo_wr_block = 0;
    assign fifo_intf_833.finish = finish;
    csv_file_dump fifo_csv_dumper_833;
    csv_file_dump cstatus_csv_dumper_833;
    df_fifo_monitor fifo_monitor_833;
    df_fifo_intf fifo_intf_834(clock,reset);
    assign fifo_intf_834.rd_en = AESL_inst_myproject.layer2_out_833_U.if_read & AESL_inst_myproject.layer2_out_833_U.if_empty_n;
    assign fifo_intf_834.wr_en = AESL_inst_myproject.layer2_out_833_U.if_write & AESL_inst_myproject.layer2_out_833_U.if_full_n;
    assign fifo_intf_834.fifo_rd_block = 0;
    assign fifo_intf_834.fifo_wr_block = 0;
    assign fifo_intf_834.finish = finish;
    csv_file_dump fifo_csv_dumper_834;
    csv_file_dump cstatus_csv_dumper_834;
    df_fifo_monitor fifo_monitor_834;
    df_fifo_intf fifo_intf_835(clock,reset);
    assign fifo_intf_835.rd_en = AESL_inst_myproject.layer2_out_834_U.if_read & AESL_inst_myproject.layer2_out_834_U.if_empty_n;
    assign fifo_intf_835.wr_en = AESL_inst_myproject.layer2_out_834_U.if_write & AESL_inst_myproject.layer2_out_834_U.if_full_n;
    assign fifo_intf_835.fifo_rd_block = 0;
    assign fifo_intf_835.fifo_wr_block = 0;
    assign fifo_intf_835.finish = finish;
    csv_file_dump fifo_csv_dumper_835;
    csv_file_dump cstatus_csv_dumper_835;
    df_fifo_monitor fifo_monitor_835;
    df_fifo_intf fifo_intf_836(clock,reset);
    assign fifo_intf_836.rd_en = AESL_inst_myproject.layer2_out_835_U.if_read & AESL_inst_myproject.layer2_out_835_U.if_empty_n;
    assign fifo_intf_836.wr_en = AESL_inst_myproject.layer2_out_835_U.if_write & AESL_inst_myproject.layer2_out_835_U.if_full_n;
    assign fifo_intf_836.fifo_rd_block = 0;
    assign fifo_intf_836.fifo_wr_block = 0;
    assign fifo_intf_836.finish = finish;
    csv_file_dump fifo_csv_dumper_836;
    csv_file_dump cstatus_csv_dumper_836;
    df_fifo_monitor fifo_monitor_836;
    df_fifo_intf fifo_intf_837(clock,reset);
    assign fifo_intf_837.rd_en = AESL_inst_myproject.layer2_out_836_U.if_read & AESL_inst_myproject.layer2_out_836_U.if_empty_n;
    assign fifo_intf_837.wr_en = AESL_inst_myproject.layer2_out_836_U.if_write & AESL_inst_myproject.layer2_out_836_U.if_full_n;
    assign fifo_intf_837.fifo_rd_block = 0;
    assign fifo_intf_837.fifo_wr_block = 0;
    assign fifo_intf_837.finish = finish;
    csv_file_dump fifo_csv_dumper_837;
    csv_file_dump cstatus_csv_dumper_837;
    df_fifo_monitor fifo_monitor_837;
    df_fifo_intf fifo_intf_838(clock,reset);
    assign fifo_intf_838.rd_en = AESL_inst_myproject.layer2_out_837_U.if_read & AESL_inst_myproject.layer2_out_837_U.if_empty_n;
    assign fifo_intf_838.wr_en = AESL_inst_myproject.layer2_out_837_U.if_write & AESL_inst_myproject.layer2_out_837_U.if_full_n;
    assign fifo_intf_838.fifo_rd_block = 0;
    assign fifo_intf_838.fifo_wr_block = 0;
    assign fifo_intf_838.finish = finish;
    csv_file_dump fifo_csv_dumper_838;
    csv_file_dump cstatus_csv_dumper_838;
    df_fifo_monitor fifo_monitor_838;
    df_fifo_intf fifo_intf_839(clock,reset);
    assign fifo_intf_839.rd_en = AESL_inst_myproject.layer2_out_838_U.if_read & AESL_inst_myproject.layer2_out_838_U.if_empty_n;
    assign fifo_intf_839.wr_en = AESL_inst_myproject.layer2_out_838_U.if_write & AESL_inst_myproject.layer2_out_838_U.if_full_n;
    assign fifo_intf_839.fifo_rd_block = 0;
    assign fifo_intf_839.fifo_wr_block = 0;
    assign fifo_intf_839.finish = finish;
    csv_file_dump fifo_csv_dumper_839;
    csv_file_dump cstatus_csv_dumper_839;
    df_fifo_monitor fifo_monitor_839;
    df_fifo_intf fifo_intf_840(clock,reset);
    assign fifo_intf_840.rd_en = AESL_inst_myproject.layer2_out_839_U.if_read & AESL_inst_myproject.layer2_out_839_U.if_empty_n;
    assign fifo_intf_840.wr_en = AESL_inst_myproject.layer2_out_839_U.if_write & AESL_inst_myproject.layer2_out_839_U.if_full_n;
    assign fifo_intf_840.fifo_rd_block = 0;
    assign fifo_intf_840.fifo_wr_block = 0;
    assign fifo_intf_840.finish = finish;
    csv_file_dump fifo_csv_dumper_840;
    csv_file_dump cstatus_csv_dumper_840;
    df_fifo_monitor fifo_monitor_840;
    df_fifo_intf fifo_intf_841(clock,reset);
    assign fifo_intf_841.rd_en = AESL_inst_myproject.layer2_out_840_U.if_read & AESL_inst_myproject.layer2_out_840_U.if_empty_n;
    assign fifo_intf_841.wr_en = AESL_inst_myproject.layer2_out_840_U.if_write & AESL_inst_myproject.layer2_out_840_U.if_full_n;
    assign fifo_intf_841.fifo_rd_block = 0;
    assign fifo_intf_841.fifo_wr_block = 0;
    assign fifo_intf_841.finish = finish;
    csv_file_dump fifo_csv_dumper_841;
    csv_file_dump cstatus_csv_dumper_841;
    df_fifo_monitor fifo_monitor_841;
    df_fifo_intf fifo_intf_842(clock,reset);
    assign fifo_intf_842.rd_en = AESL_inst_myproject.layer2_out_841_U.if_read & AESL_inst_myproject.layer2_out_841_U.if_empty_n;
    assign fifo_intf_842.wr_en = AESL_inst_myproject.layer2_out_841_U.if_write & AESL_inst_myproject.layer2_out_841_U.if_full_n;
    assign fifo_intf_842.fifo_rd_block = 0;
    assign fifo_intf_842.fifo_wr_block = 0;
    assign fifo_intf_842.finish = finish;
    csv_file_dump fifo_csv_dumper_842;
    csv_file_dump cstatus_csv_dumper_842;
    df_fifo_monitor fifo_monitor_842;
    df_fifo_intf fifo_intf_843(clock,reset);
    assign fifo_intf_843.rd_en = AESL_inst_myproject.layer2_out_842_U.if_read & AESL_inst_myproject.layer2_out_842_U.if_empty_n;
    assign fifo_intf_843.wr_en = AESL_inst_myproject.layer2_out_842_U.if_write & AESL_inst_myproject.layer2_out_842_U.if_full_n;
    assign fifo_intf_843.fifo_rd_block = 0;
    assign fifo_intf_843.fifo_wr_block = 0;
    assign fifo_intf_843.finish = finish;
    csv_file_dump fifo_csv_dumper_843;
    csv_file_dump cstatus_csv_dumper_843;
    df_fifo_monitor fifo_monitor_843;
    df_fifo_intf fifo_intf_844(clock,reset);
    assign fifo_intf_844.rd_en = AESL_inst_myproject.layer2_out_843_U.if_read & AESL_inst_myproject.layer2_out_843_U.if_empty_n;
    assign fifo_intf_844.wr_en = AESL_inst_myproject.layer2_out_843_U.if_write & AESL_inst_myproject.layer2_out_843_U.if_full_n;
    assign fifo_intf_844.fifo_rd_block = 0;
    assign fifo_intf_844.fifo_wr_block = 0;
    assign fifo_intf_844.finish = finish;
    csv_file_dump fifo_csv_dumper_844;
    csv_file_dump cstatus_csv_dumper_844;
    df_fifo_monitor fifo_monitor_844;
    df_fifo_intf fifo_intf_845(clock,reset);
    assign fifo_intf_845.rd_en = AESL_inst_myproject.layer2_out_844_U.if_read & AESL_inst_myproject.layer2_out_844_U.if_empty_n;
    assign fifo_intf_845.wr_en = AESL_inst_myproject.layer2_out_844_U.if_write & AESL_inst_myproject.layer2_out_844_U.if_full_n;
    assign fifo_intf_845.fifo_rd_block = 0;
    assign fifo_intf_845.fifo_wr_block = 0;
    assign fifo_intf_845.finish = finish;
    csv_file_dump fifo_csv_dumper_845;
    csv_file_dump cstatus_csv_dumper_845;
    df_fifo_monitor fifo_monitor_845;
    df_fifo_intf fifo_intf_846(clock,reset);
    assign fifo_intf_846.rd_en = AESL_inst_myproject.layer2_out_845_U.if_read & AESL_inst_myproject.layer2_out_845_U.if_empty_n;
    assign fifo_intf_846.wr_en = AESL_inst_myproject.layer2_out_845_U.if_write & AESL_inst_myproject.layer2_out_845_U.if_full_n;
    assign fifo_intf_846.fifo_rd_block = 0;
    assign fifo_intf_846.fifo_wr_block = 0;
    assign fifo_intf_846.finish = finish;
    csv_file_dump fifo_csv_dumper_846;
    csv_file_dump cstatus_csv_dumper_846;
    df_fifo_monitor fifo_monitor_846;
    df_fifo_intf fifo_intf_847(clock,reset);
    assign fifo_intf_847.rd_en = AESL_inst_myproject.layer2_out_846_U.if_read & AESL_inst_myproject.layer2_out_846_U.if_empty_n;
    assign fifo_intf_847.wr_en = AESL_inst_myproject.layer2_out_846_U.if_write & AESL_inst_myproject.layer2_out_846_U.if_full_n;
    assign fifo_intf_847.fifo_rd_block = 0;
    assign fifo_intf_847.fifo_wr_block = 0;
    assign fifo_intf_847.finish = finish;
    csv_file_dump fifo_csv_dumper_847;
    csv_file_dump cstatus_csv_dumper_847;
    df_fifo_monitor fifo_monitor_847;
    df_fifo_intf fifo_intf_848(clock,reset);
    assign fifo_intf_848.rd_en = AESL_inst_myproject.layer2_out_847_U.if_read & AESL_inst_myproject.layer2_out_847_U.if_empty_n;
    assign fifo_intf_848.wr_en = AESL_inst_myproject.layer2_out_847_U.if_write & AESL_inst_myproject.layer2_out_847_U.if_full_n;
    assign fifo_intf_848.fifo_rd_block = 0;
    assign fifo_intf_848.fifo_wr_block = 0;
    assign fifo_intf_848.finish = finish;
    csv_file_dump fifo_csv_dumper_848;
    csv_file_dump cstatus_csv_dumper_848;
    df_fifo_monitor fifo_monitor_848;
    df_fifo_intf fifo_intf_849(clock,reset);
    assign fifo_intf_849.rd_en = AESL_inst_myproject.layer2_out_848_U.if_read & AESL_inst_myproject.layer2_out_848_U.if_empty_n;
    assign fifo_intf_849.wr_en = AESL_inst_myproject.layer2_out_848_U.if_write & AESL_inst_myproject.layer2_out_848_U.if_full_n;
    assign fifo_intf_849.fifo_rd_block = 0;
    assign fifo_intf_849.fifo_wr_block = 0;
    assign fifo_intf_849.finish = finish;
    csv_file_dump fifo_csv_dumper_849;
    csv_file_dump cstatus_csv_dumper_849;
    df_fifo_monitor fifo_monitor_849;
    df_fifo_intf fifo_intf_850(clock,reset);
    assign fifo_intf_850.rd_en = AESL_inst_myproject.layer2_out_849_U.if_read & AESL_inst_myproject.layer2_out_849_U.if_empty_n;
    assign fifo_intf_850.wr_en = AESL_inst_myproject.layer2_out_849_U.if_write & AESL_inst_myproject.layer2_out_849_U.if_full_n;
    assign fifo_intf_850.fifo_rd_block = 0;
    assign fifo_intf_850.fifo_wr_block = 0;
    assign fifo_intf_850.finish = finish;
    csv_file_dump fifo_csv_dumper_850;
    csv_file_dump cstatus_csv_dumper_850;
    df_fifo_monitor fifo_monitor_850;
    df_fifo_intf fifo_intf_851(clock,reset);
    assign fifo_intf_851.rd_en = AESL_inst_myproject.layer2_out_850_U.if_read & AESL_inst_myproject.layer2_out_850_U.if_empty_n;
    assign fifo_intf_851.wr_en = AESL_inst_myproject.layer2_out_850_U.if_write & AESL_inst_myproject.layer2_out_850_U.if_full_n;
    assign fifo_intf_851.fifo_rd_block = 0;
    assign fifo_intf_851.fifo_wr_block = 0;
    assign fifo_intf_851.finish = finish;
    csv_file_dump fifo_csv_dumper_851;
    csv_file_dump cstatus_csv_dumper_851;
    df_fifo_monitor fifo_monitor_851;
    df_fifo_intf fifo_intf_852(clock,reset);
    assign fifo_intf_852.rd_en = AESL_inst_myproject.layer2_out_851_U.if_read & AESL_inst_myproject.layer2_out_851_U.if_empty_n;
    assign fifo_intf_852.wr_en = AESL_inst_myproject.layer2_out_851_U.if_write & AESL_inst_myproject.layer2_out_851_U.if_full_n;
    assign fifo_intf_852.fifo_rd_block = 0;
    assign fifo_intf_852.fifo_wr_block = 0;
    assign fifo_intf_852.finish = finish;
    csv_file_dump fifo_csv_dumper_852;
    csv_file_dump cstatus_csv_dumper_852;
    df_fifo_monitor fifo_monitor_852;
    df_fifo_intf fifo_intf_853(clock,reset);
    assign fifo_intf_853.rd_en = AESL_inst_myproject.layer2_out_852_U.if_read & AESL_inst_myproject.layer2_out_852_U.if_empty_n;
    assign fifo_intf_853.wr_en = AESL_inst_myproject.layer2_out_852_U.if_write & AESL_inst_myproject.layer2_out_852_U.if_full_n;
    assign fifo_intf_853.fifo_rd_block = 0;
    assign fifo_intf_853.fifo_wr_block = 0;
    assign fifo_intf_853.finish = finish;
    csv_file_dump fifo_csv_dumper_853;
    csv_file_dump cstatus_csv_dumper_853;
    df_fifo_monitor fifo_monitor_853;
    df_fifo_intf fifo_intf_854(clock,reset);
    assign fifo_intf_854.rd_en = AESL_inst_myproject.layer2_out_853_U.if_read & AESL_inst_myproject.layer2_out_853_U.if_empty_n;
    assign fifo_intf_854.wr_en = AESL_inst_myproject.layer2_out_853_U.if_write & AESL_inst_myproject.layer2_out_853_U.if_full_n;
    assign fifo_intf_854.fifo_rd_block = 0;
    assign fifo_intf_854.fifo_wr_block = 0;
    assign fifo_intf_854.finish = finish;
    csv_file_dump fifo_csv_dumper_854;
    csv_file_dump cstatus_csv_dumper_854;
    df_fifo_monitor fifo_monitor_854;
    df_fifo_intf fifo_intf_855(clock,reset);
    assign fifo_intf_855.rd_en = AESL_inst_myproject.layer2_out_854_U.if_read & AESL_inst_myproject.layer2_out_854_U.if_empty_n;
    assign fifo_intf_855.wr_en = AESL_inst_myproject.layer2_out_854_U.if_write & AESL_inst_myproject.layer2_out_854_U.if_full_n;
    assign fifo_intf_855.fifo_rd_block = 0;
    assign fifo_intf_855.fifo_wr_block = 0;
    assign fifo_intf_855.finish = finish;
    csv_file_dump fifo_csv_dumper_855;
    csv_file_dump cstatus_csv_dumper_855;
    df_fifo_monitor fifo_monitor_855;
    df_fifo_intf fifo_intf_856(clock,reset);
    assign fifo_intf_856.rd_en = AESL_inst_myproject.layer2_out_855_U.if_read & AESL_inst_myproject.layer2_out_855_U.if_empty_n;
    assign fifo_intf_856.wr_en = AESL_inst_myproject.layer2_out_855_U.if_write & AESL_inst_myproject.layer2_out_855_U.if_full_n;
    assign fifo_intf_856.fifo_rd_block = 0;
    assign fifo_intf_856.fifo_wr_block = 0;
    assign fifo_intf_856.finish = finish;
    csv_file_dump fifo_csv_dumper_856;
    csv_file_dump cstatus_csv_dumper_856;
    df_fifo_monitor fifo_monitor_856;
    df_fifo_intf fifo_intf_857(clock,reset);
    assign fifo_intf_857.rd_en = AESL_inst_myproject.layer2_out_856_U.if_read & AESL_inst_myproject.layer2_out_856_U.if_empty_n;
    assign fifo_intf_857.wr_en = AESL_inst_myproject.layer2_out_856_U.if_write & AESL_inst_myproject.layer2_out_856_U.if_full_n;
    assign fifo_intf_857.fifo_rd_block = 0;
    assign fifo_intf_857.fifo_wr_block = 0;
    assign fifo_intf_857.finish = finish;
    csv_file_dump fifo_csv_dumper_857;
    csv_file_dump cstatus_csv_dumper_857;
    df_fifo_monitor fifo_monitor_857;
    df_fifo_intf fifo_intf_858(clock,reset);
    assign fifo_intf_858.rd_en = AESL_inst_myproject.layer2_out_857_U.if_read & AESL_inst_myproject.layer2_out_857_U.if_empty_n;
    assign fifo_intf_858.wr_en = AESL_inst_myproject.layer2_out_857_U.if_write & AESL_inst_myproject.layer2_out_857_U.if_full_n;
    assign fifo_intf_858.fifo_rd_block = 0;
    assign fifo_intf_858.fifo_wr_block = 0;
    assign fifo_intf_858.finish = finish;
    csv_file_dump fifo_csv_dumper_858;
    csv_file_dump cstatus_csv_dumper_858;
    df_fifo_monitor fifo_monitor_858;
    df_fifo_intf fifo_intf_859(clock,reset);
    assign fifo_intf_859.rd_en = AESL_inst_myproject.layer2_out_858_U.if_read & AESL_inst_myproject.layer2_out_858_U.if_empty_n;
    assign fifo_intf_859.wr_en = AESL_inst_myproject.layer2_out_858_U.if_write & AESL_inst_myproject.layer2_out_858_U.if_full_n;
    assign fifo_intf_859.fifo_rd_block = 0;
    assign fifo_intf_859.fifo_wr_block = 0;
    assign fifo_intf_859.finish = finish;
    csv_file_dump fifo_csv_dumper_859;
    csv_file_dump cstatus_csv_dumper_859;
    df_fifo_monitor fifo_monitor_859;
    df_fifo_intf fifo_intf_860(clock,reset);
    assign fifo_intf_860.rd_en = AESL_inst_myproject.layer2_out_859_U.if_read & AESL_inst_myproject.layer2_out_859_U.if_empty_n;
    assign fifo_intf_860.wr_en = AESL_inst_myproject.layer2_out_859_U.if_write & AESL_inst_myproject.layer2_out_859_U.if_full_n;
    assign fifo_intf_860.fifo_rd_block = 0;
    assign fifo_intf_860.fifo_wr_block = 0;
    assign fifo_intf_860.finish = finish;
    csv_file_dump fifo_csv_dumper_860;
    csv_file_dump cstatus_csv_dumper_860;
    df_fifo_monitor fifo_monitor_860;
    df_fifo_intf fifo_intf_861(clock,reset);
    assign fifo_intf_861.rd_en = AESL_inst_myproject.layer2_out_860_U.if_read & AESL_inst_myproject.layer2_out_860_U.if_empty_n;
    assign fifo_intf_861.wr_en = AESL_inst_myproject.layer2_out_860_U.if_write & AESL_inst_myproject.layer2_out_860_U.if_full_n;
    assign fifo_intf_861.fifo_rd_block = 0;
    assign fifo_intf_861.fifo_wr_block = 0;
    assign fifo_intf_861.finish = finish;
    csv_file_dump fifo_csv_dumper_861;
    csv_file_dump cstatus_csv_dumper_861;
    df_fifo_monitor fifo_monitor_861;
    df_fifo_intf fifo_intf_862(clock,reset);
    assign fifo_intf_862.rd_en = AESL_inst_myproject.layer2_out_861_U.if_read & AESL_inst_myproject.layer2_out_861_U.if_empty_n;
    assign fifo_intf_862.wr_en = AESL_inst_myproject.layer2_out_861_U.if_write & AESL_inst_myproject.layer2_out_861_U.if_full_n;
    assign fifo_intf_862.fifo_rd_block = 0;
    assign fifo_intf_862.fifo_wr_block = 0;
    assign fifo_intf_862.finish = finish;
    csv_file_dump fifo_csv_dumper_862;
    csv_file_dump cstatus_csv_dumper_862;
    df_fifo_monitor fifo_monitor_862;
    df_fifo_intf fifo_intf_863(clock,reset);
    assign fifo_intf_863.rd_en = AESL_inst_myproject.layer2_out_862_U.if_read & AESL_inst_myproject.layer2_out_862_U.if_empty_n;
    assign fifo_intf_863.wr_en = AESL_inst_myproject.layer2_out_862_U.if_write & AESL_inst_myproject.layer2_out_862_U.if_full_n;
    assign fifo_intf_863.fifo_rd_block = 0;
    assign fifo_intf_863.fifo_wr_block = 0;
    assign fifo_intf_863.finish = finish;
    csv_file_dump fifo_csv_dumper_863;
    csv_file_dump cstatus_csv_dumper_863;
    df_fifo_monitor fifo_monitor_863;
    df_fifo_intf fifo_intf_864(clock,reset);
    assign fifo_intf_864.rd_en = AESL_inst_myproject.layer2_out_863_U.if_read & AESL_inst_myproject.layer2_out_863_U.if_empty_n;
    assign fifo_intf_864.wr_en = AESL_inst_myproject.layer2_out_863_U.if_write & AESL_inst_myproject.layer2_out_863_U.if_full_n;
    assign fifo_intf_864.fifo_rd_block = 0;
    assign fifo_intf_864.fifo_wr_block = 0;
    assign fifo_intf_864.finish = finish;
    csv_file_dump fifo_csv_dumper_864;
    csv_file_dump cstatus_csv_dumper_864;
    df_fifo_monitor fifo_monitor_864;
    df_fifo_intf fifo_intf_865(clock,reset);
    assign fifo_intf_865.rd_en = AESL_inst_myproject.layer2_out_864_U.if_read & AESL_inst_myproject.layer2_out_864_U.if_empty_n;
    assign fifo_intf_865.wr_en = AESL_inst_myproject.layer2_out_864_U.if_write & AESL_inst_myproject.layer2_out_864_U.if_full_n;
    assign fifo_intf_865.fifo_rd_block = 0;
    assign fifo_intf_865.fifo_wr_block = 0;
    assign fifo_intf_865.finish = finish;
    csv_file_dump fifo_csv_dumper_865;
    csv_file_dump cstatus_csv_dumper_865;
    df_fifo_monitor fifo_monitor_865;
    df_fifo_intf fifo_intf_866(clock,reset);
    assign fifo_intf_866.rd_en = AESL_inst_myproject.layer2_out_865_U.if_read & AESL_inst_myproject.layer2_out_865_U.if_empty_n;
    assign fifo_intf_866.wr_en = AESL_inst_myproject.layer2_out_865_U.if_write & AESL_inst_myproject.layer2_out_865_U.if_full_n;
    assign fifo_intf_866.fifo_rd_block = 0;
    assign fifo_intf_866.fifo_wr_block = 0;
    assign fifo_intf_866.finish = finish;
    csv_file_dump fifo_csv_dumper_866;
    csv_file_dump cstatus_csv_dumper_866;
    df_fifo_monitor fifo_monitor_866;
    df_fifo_intf fifo_intf_867(clock,reset);
    assign fifo_intf_867.rd_en = AESL_inst_myproject.layer2_out_866_U.if_read & AESL_inst_myproject.layer2_out_866_U.if_empty_n;
    assign fifo_intf_867.wr_en = AESL_inst_myproject.layer2_out_866_U.if_write & AESL_inst_myproject.layer2_out_866_U.if_full_n;
    assign fifo_intf_867.fifo_rd_block = 0;
    assign fifo_intf_867.fifo_wr_block = 0;
    assign fifo_intf_867.finish = finish;
    csv_file_dump fifo_csv_dumper_867;
    csv_file_dump cstatus_csv_dumper_867;
    df_fifo_monitor fifo_monitor_867;
    df_fifo_intf fifo_intf_868(clock,reset);
    assign fifo_intf_868.rd_en = AESL_inst_myproject.layer2_out_867_U.if_read & AESL_inst_myproject.layer2_out_867_U.if_empty_n;
    assign fifo_intf_868.wr_en = AESL_inst_myproject.layer2_out_867_U.if_write & AESL_inst_myproject.layer2_out_867_U.if_full_n;
    assign fifo_intf_868.fifo_rd_block = 0;
    assign fifo_intf_868.fifo_wr_block = 0;
    assign fifo_intf_868.finish = finish;
    csv_file_dump fifo_csv_dumper_868;
    csv_file_dump cstatus_csv_dumper_868;
    df_fifo_monitor fifo_monitor_868;
    df_fifo_intf fifo_intf_869(clock,reset);
    assign fifo_intf_869.rd_en = AESL_inst_myproject.layer2_out_868_U.if_read & AESL_inst_myproject.layer2_out_868_U.if_empty_n;
    assign fifo_intf_869.wr_en = AESL_inst_myproject.layer2_out_868_U.if_write & AESL_inst_myproject.layer2_out_868_U.if_full_n;
    assign fifo_intf_869.fifo_rd_block = 0;
    assign fifo_intf_869.fifo_wr_block = 0;
    assign fifo_intf_869.finish = finish;
    csv_file_dump fifo_csv_dumper_869;
    csv_file_dump cstatus_csv_dumper_869;
    df_fifo_monitor fifo_monitor_869;
    df_fifo_intf fifo_intf_870(clock,reset);
    assign fifo_intf_870.rd_en = AESL_inst_myproject.layer2_out_869_U.if_read & AESL_inst_myproject.layer2_out_869_U.if_empty_n;
    assign fifo_intf_870.wr_en = AESL_inst_myproject.layer2_out_869_U.if_write & AESL_inst_myproject.layer2_out_869_U.if_full_n;
    assign fifo_intf_870.fifo_rd_block = 0;
    assign fifo_intf_870.fifo_wr_block = 0;
    assign fifo_intf_870.finish = finish;
    csv_file_dump fifo_csv_dumper_870;
    csv_file_dump cstatus_csv_dumper_870;
    df_fifo_monitor fifo_monitor_870;
    df_fifo_intf fifo_intf_871(clock,reset);
    assign fifo_intf_871.rd_en = AESL_inst_myproject.layer2_out_870_U.if_read & AESL_inst_myproject.layer2_out_870_U.if_empty_n;
    assign fifo_intf_871.wr_en = AESL_inst_myproject.layer2_out_870_U.if_write & AESL_inst_myproject.layer2_out_870_U.if_full_n;
    assign fifo_intf_871.fifo_rd_block = 0;
    assign fifo_intf_871.fifo_wr_block = 0;
    assign fifo_intf_871.finish = finish;
    csv_file_dump fifo_csv_dumper_871;
    csv_file_dump cstatus_csv_dumper_871;
    df_fifo_monitor fifo_monitor_871;
    df_fifo_intf fifo_intf_872(clock,reset);
    assign fifo_intf_872.rd_en = AESL_inst_myproject.layer2_out_871_U.if_read & AESL_inst_myproject.layer2_out_871_U.if_empty_n;
    assign fifo_intf_872.wr_en = AESL_inst_myproject.layer2_out_871_U.if_write & AESL_inst_myproject.layer2_out_871_U.if_full_n;
    assign fifo_intf_872.fifo_rd_block = 0;
    assign fifo_intf_872.fifo_wr_block = 0;
    assign fifo_intf_872.finish = finish;
    csv_file_dump fifo_csv_dumper_872;
    csv_file_dump cstatus_csv_dumper_872;
    df_fifo_monitor fifo_monitor_872;
    df_fifo_intf fifo_intf_873(clock,reset);
    assign fifo_intf_873.rd_en = AESL_inst_myproject.layer2_out_872_U.if_read & AESL_inst_myproject.layer2_out_872_U.if_empty_n;
    assign fifo_intf_873.wr_en = AESL_inst_myproject.layer2_out_872_U.if_write & AESL_inst_myproject.layer2_out_872_U.if_full_n;
    assign fifo_intf_873.fifo_rd_block = 0;
    assign fifo_intf_873.fifo_wr_block = 0;
    assign fifo_intf_873.finish = finish;
    csv_file_dump fifo_csv_dumper_873;
    csv_file_dump cstatus_csv_dumper_873;
    df_fifo_monitor fifo_monitor_873;
    df_fifo_intf fifo_intf_874(clock,reset);
    assign fifo_intf_874.rd_en = AESL_inst_myproject.layer2_out_873_U.if_read & AESL_inst_myproject.layer2_out_873_U.if_empty_n;
    assign fifo_intf_874.wr_en = AESL_inst_myproject.layer2_out_873_U.if_write & AESL_inst_myproject.layer2_out_873_U.if_full_n;
    assign fifo_intf_874.fifo_rd_block = 0;
    assign fifo_intf_874.fifo_wr_block = 0;
    assign fifo_intf_874.finish = finish;
    csv_file_dump fifo_csv_dumper_874;
    csv_file_dump cstatus_csv_dumper_874;
    df_fifo_monitor fifo_monitor_874;
    df_fifo_intf fifo_intf_875(clock,reset);
    assign fifo_intf_875.rd_en = AESL_inst_myproject.layer2_out_874_U.if_read & AESL_inst_myproject.layer2_out_874_U.if_empty_n;
    assign fifo_intf_875.wr_en = AESL_inst_myproject.layer2_out_874_U.if_write & AESL_inst_myproject.layer2_out_874_U.if_full_n;
    assign fifo_intf_875.fifo_rd_block = 0;
    assign fifo_intf_875.fifo_wr_block = 0;
    assign fifo_intf_875.finish = finish;
    csv_file_dump fifo_csv_dumper_875;
    csv_file_dump cstatus_csv_dumper_875;
    df_fifo_monitor fifo_monitor_875;
    df_fifo_intf fifo_intf_876(clock,reset);
    assign fifo_intf_876.rd_en = AESL_inst_myproject.layer2_out_875_U.if_read & AESL_inst_myproject.layer2_out_875_U.if_empty_n;
    assign fifo_intf_876.wr_en = AESL_inst_myproject.layer2_out_875_U.if_write & AESL_inst_myproject.layer2_out_875_U.if_full_n;
    assign fifo_intf_876.fifo_rd_block = 0;
    assign fifo_intf_876.fifo_wr_block = 0;
    assign fifo_intf_876.finish = finish;
    csv_file_dump fifo_csv_dumper_876;
    csv_file_dump cstatus_csv_dumper_876;
    df_fifo_monitor fifo_monitor_876;
    df_fifo_intf fifo_intf_877(clock,reset);
    assign fifo_intf_877.rd_en = AESL_inst_myproject.layer2_out_876_U.if_read & AESL_inst_myproject.layer2_out_876_U.if_empty_n;
    assign fifo_intf_877.wr_en = AESL_inst_myproject.layer2_out_876_U.if_write & AESL_inst_myproject.layer2_out_876_U.if_full_n;
    assign fifo_intf_877.fifo_rd_block = 0;
    assign fifo_intf_877.fifo_wr_block = 0;
    assign fifo_intf_877.finish = finish;
    csv_file_dump fifo_csv_dumper_877;
    csv_file_dump cstatus_csv_dumper_877;
    df_fifo_monitor fifo_monitor_877;
    df_fifo_intf fifo_intf_878(clock,reset);
    assign fifo_intf_878.rd_en = AESL_inst_myproject.layer2_out_877_U.if_read & AESL_inst_myproject.layer2_out_877_U.if_empty_n;
    assign fifo_intf_878.wr_en = AESL_inst_myproject.layer2_out_877_U.if_write & AESL_inst_myproject.layer2_out_877_U.if_full_n;
    assign fifo_intf_878.fifo_rd_block = 0;
    assign fifo_intf_878.fifo_wr_block = 0;
    assign fifo_intf_878.finish = finish;
    csv_file_dump fifo_csv_dumper_878;
    csv_file_dump cstatus_csv_dumper_878;
    df_fifo_monitor fifo_monitor_878;
    df_fifo_intf fifo_intf_879(clock,reset);
    assign fifo_intf_879.rd_en = AESL_inst_myproject.layer2_out_878_U.if_read & AESL_inst_myproject.layer2_out_878_U.if_empty_n;
    assign fifo_intf_879.wr_en = AESL_inst_myproject.layer2_out_878_U.if_write & AESL_inst_myproject.layer2_out_878_U.if_full_n;
    assign fifo_intf_879.fifo_rd_block = 0;
    assign fifo_intf_879.fifo_wr_block = 0;
    assign fifo_intf_879.finish = finish;
    csv_file_dump fifo_csv_dumper_879;
    csv_file_dump cstatus_csv_dumper_879;
    df_fifo_monitor fifo_monitor_879;
    df_fifo_intf fifo_intf_880(clock,reset);
    assign fifo_intf_880.rd_en = AESL_inst_myproject.layer2_out_879_U.if_read & AESL_inst_myproject.layer2_out_879_U.if_empty_n;
    assign fifo_intf_880.wr_en = AESL_inst_myproject.layer2_out_879_U.if_write & AESL_inst_myproject.layer2_out_879_U.if_full_n;
    assign fifo_intf_880.fifo_rd_block = 0;
    assign fifo_intf_880.fifo_wr_block = 0;
    assign fifo_intf_880.finish = finish;
    csv_file_dump fifo_csv_dumper_880;
    csv_file_dump cstatus_csv_dumper_880;
    df_fifo_monitor fifo_monitor_880;
    df_fifo_intf fifo_intf_881(clock,reset);
    assign fifo_intf_881.rd_en = AESL_inst_myproject.layer2_out_880_U.if_read & AESL_inst_myproject.layer2_out_880_U.if_empty_n;
    assign fifo_intf_881.wr_en = AESL_inst_myproject.layer2_out_880_U.if_write & AESL_inst_myproject.layer2_out_880_U.if_full_n;
    assign fifo_intf_881.fifo_rd_block = 0;
    assign fifo_intf_881.fifo_wr_block = 0;
    assign fifo_intf_881.finish = finish;
    csv_file_dump fifo_csv_dumper_881;
    csv_file_dump cstatus_csv_dumper_881;
    df_fifo_monitor fifo_monitor_881;
    df_fifo_intf fifo_intf_882(clock,reset);
    assign fifo_intf_882.rd_en = AESL_inst_myproject.layer2_out_881_U.if_read & AESL_inst_myproject.layer2_out_881_U.if_empty_n;
    assign fifo_intf_882.wr_en = AESL_inst_myproject.layer2_out_881_U.if_write & AESL_inst_myproject.layer2_out_881_U.if_full_n;
    assign fifo_intf_882.fifo_rd_block = 0;
    assign fifo_intf_882.fifo_wr_block = 0;
    assign fifo_intf_882.finish = finish;
    csv_file_dump fifo_csv_dumper_882;
    csv_file_dump cstatus_csv_dumper_882;
    df_fifo_monitor fifo_monitor_882;
    df_fifo_intf fifo_intf_883(clock,reset);
    assign fifo_intf_883.rd_en = AESL_inst_myproject.layer2_out_882_U.if_read & AESL_inst_myproject.layer2_out_882_U.if_empty_n;
    assign fifo_intf_883.wr_en = AESL_inst_myproject.layer2_out_882_U.if_write & AESL_inst_myproject.layer2_out_882_U.if_full_n;
    assign fifo_intf_883.fifo_rd_block = 0;
    assign fifo_intf_883.fifo_wr_block = 0;
    assign fifo_intf_883.finish = finish;
    csv_file_dump fifo_csv_dumper_883;
    csv_file_dump cstatus_csv_dumper_883;
    df_fifo_monitor fifo_monitor_883;
    df_fifo_intf fifo_intf_884(clock,reset);
    assign fifo_intf_884.rd_en = AESL_inst_myproject.layer2_out_883_U.if_read & AESL_inst_myproject.layer2_out_883_U.if_empty_n;
    assign fifo_intf_884.wr_en = AESL_inst_myproject.layer2_out_883_U.if_write & AESL_inst_myproject.layer2_out_883_U.if_full_n;
    assign fifo_intf_884.fifo_rd_block = 0;
    assign fifo_intf_884.fifo_wr_block = 0;
    assign fifo_intf_884.finish = finish;
    csv_file_dump fifo_csv_dumper_884;
    csv_file_dump cstatus_csv_dumper_884;
    df_fifo_monitor fifo_monitor_884;
    df_fifo_intf fifo_intf_885(clock,reset);
    assign fifo_intf_885.rd_en = AESL_inst_myproject.layer2_out_884_U.if_read & AESL_inst_myproject.layer2_out_884_U.if_empty_n;
    assign fifo_intf_885.wr_en = AESL_inst_myproject.layer2_out_884_U.if_write & AESL_inst_myproject.layer2_out_884_U.if_full_n;
    assign fifo_intf_885.fifo_rd_block = 0;
    assign fifo_intf_885.fifo_wr_block = 0;
    assign fifo_intf_885.finish = finish;
    csv_file_dump fifo_csv_dumper_885;
    csv_file_dump cstatus_csv_dumper_885;
    df_fifo_monitor fifo_monitor_885;
    df_fifo_intf fifo_intf_886(clock,reset);
    assign fifo_intf_886.rd_en = AESL_inst_myproject.layer2_out_885_U.if_read & AESL_inst_myproject.layer2_out_885_U.if_empty_n;
    assign fifo_intf_886.wr_en = AESL_inst_myproject.layer2_out_885_U.if_write & AESL_inst_myproject.layer2_out_885_U.if_full_n;
    assign fifo_intf_886.fifo_rd_block = 0;
    assign fifo_intf_886.fifo_wr_block = 0;
    assign fifo_intf_886.finish = finish;
    csv_file_dump fifo_csv_dumper_886;
    csv_file_dump cstatus_csv_dumper_886;
    df_fifo_monitor fifo_monitor_886;
    df_fifo_intf fifo_intf_887(clock,reset);
    assign fifo_intf_887.rd_en = AESL_inst_myproject.layer2_out_886_U.if_read & AESL_inst_myproject.layer2_out_886_U.if_empty_n;
    assign fifo_intf_887.wr_en = AESL_inst_myproject.layer2_out_886_U.if_write & AESL_inst_myproject.layer2_out_886_U.if_full_n;
    assign fifo_intf_887.fifo_rd_block = 0;
    assign fifo_intf_887.fifo_wr_block = 0;
    assign fifo_intf_887.finish = finish;
    csv_file_dump fifo_csv_dumper_887;
    csv_file_dump cstatus_csv_dumper_887;
    df_fifo_monitor fifo_monitor_887;
    df_fifo_intf fifo_intf_888(clock,reset);
    assign fifo_intf_888.rd_en = AESL_inst_myproject.layer2_out_887_U.if_read & AESL_inst_myproject.layer2_out_887_U.if_empty_n;
    assign fifo_intf_888.wr_en = AESL_inst_myproject.layer2_out_887_U.if_write & AESL_inst_myproject.layer2_out_887_U.if_full_n;
    assign fifo_intf_888.fifo_rd_block = 0;
    assign fifo_intf_888.fifo_wr_block = 0;
    assign fifo_intf_888.finish = finish;
    csv_file_dump fifo_csv_dumper_888;
    csv_file_dump cstatus_csv_dumper_888;
    df_fifo_monitor fifo_monitor_888;
    df_fifo_intf fifo_intf_889(clock,reset);
    assign fifo_intf_889.rd_en = AESL_inst_myproject.layer2_out_888_U.if_read & AESL_inst_myproject.layer2_out_888_U.if_empty_n;
    assign fifo_intf_889.wr_en = AESL_inst_myproject.layer2_out_888_U.if_write & AESL_inst_myproject.layer2_out_888_U.if_full_n;
    assign fifo_intf_889.fifo_rd_block = 0;
    assign fifo_intf_889.fifo_wr_block = 0;
    assign fifo_intf_889.finish = finish;
    csv_file_dump fifo_csv_dumper_889;
    csv_file_dump cstatus_csv_dumper_889;
    df_fifo_monitor fifo_monitor_889;
    df_fifo_intf fifo_intf_890(clock,reset);
    assign fifo_intf_890.rd_en = AESL_inst_myproject.layer2_out_889_U.if_read & AESL_inst_myproject.layer2_out_889_U.if_empty_n;
    assign fifo_intf_890.wr_en = AESL_inst_myproject.layer2_out_889_U.if_write & AESL_inst_myproject.layer2_out_889_U.if_full_n;
    assign fifo_intf_890.fifo_rd_block = 0;
    assign fifo_intf_890.fifo_wr_block = 0;
    assign fifo_intf_890.finish = finish;
    csv_file_dump fifo_csv_dumper_890;
    csv_file_dump cstatus_csv_dumper_890;
    df_fifo_monitor fifo_monitor_890;
    df_fifo_intf fifo_intf_891(clock,reset);
    assign fifo_intf_891.rd_en = AESL_inst_myproject.layer2_out_890_U.if_read & AESL_inst_myproject.layer2_out_890_U.if_empty_n;
    assign fifo_intf_891.wr_en = AESL_inst_myproject.layer2_out_890_U.if_write & AESL_inst_myproject.layer2_out_890_U.if_full_n;
    assign fifo_intf_891.fifo_rd_block = 0;
    assign fifo_intf_891.fifo_wr_block = 0;
    assign fifo_intf_891.finish = finish;
    csv_file_dump fifo_csv_dumper_891;
    csv_file_dump cstatus_csv_dumper_891;
    df_fifo_monitor fifo_monitor_891;
    df_fifo_intf fifo_intf_892(clock,reset);
    assign fifo_intf_892.rd_en = AESL_inst_myproject.layer2_out_891_U.if_read & AESL_inst_myproject.layer2_out_891_U.if_empty_n;
    assign fifo_intf_892.wr_en = AESL_inst_myproject.layer2_out_891_U.if_write & AESL_inst_myproject.layer2_out_891_U.if_full_n;
    assign fifo_intf_892.fifo_rd_block = 0;
    assign fifo_intf_892.fifo_wr_block = 0;
    assign fifo_intf_892.finish = finish;
    csv_file_dump fifo_csv_dumper_892;
    csv_file_dump cstatus_csv_dumper_892;
    df_fifo_monitor fifo_monitor_892;
    df_fifo_intf fifo_intf_893(clock,reset);
    assign fifo_intf_893.rd_en = AESL_inst_myproject.layer2_out_892_U.if_read & AESL_inst_myproject.layer2_out_892_U.if_empty_n;
    assign fifo_intf_893.wr_en = AESL_inst_myproject.layer2_out_892_U.if_write & AESL_inst_myproject.layer2_out_892_U.if_full_n;
    assign fifo_intf_893.fifo_rd_block = 0;
    assign fifo_intf_893.fifo_wr_block = 0;
    assign fifo_intf_893.finish = finish;
    csv_file_dump fifo_csv_dumper_893;
    csv_file_dump cstatus_csv_dumper_893;
    df_fifo_monitor fifo_monitor_893;
    df_fifo_intf fifo_intf_894(clock,reset);
    assign fifo_intf_894.rd_en = AESL_inst_myproject.layer2_out_893_U.if_read & AESL_inst_myproject.layer2_out_893_U.if_empty_n;
    assign fifo_intf_894.wr_en = AESL_inst_myproject.layer2_out_893_U.if_write & AESL_inst_myproject.layer2_out_893_U.if_full_n;
    assign fifo_intf_894.fifo_rd_block = 0;
    assign fifo_intf_894.fifo_wr_block = 0;
    assign fifo_intf_894.finish = finish;
    csv_file_dump fifo_csv_dumper_894;
    csv_file_dump cstatus_csv_dumper_894;
    df_fifo_monitor fifo_monitor_894;
    df_fifo_intf fifo_intf_895(clock,reset);
    assign fifo_intf_895.rd_en = AESL_inst_myproject.layer2_out_894_U.if_read & AESL_inst_myproject.layer2_out_894_U.if_empty_n;
    assign fifo_intf_895.wr_en = AESL_inst_myproject.layer2_out_894_U.if_write & AESL_inst_myproject.layer2_out_894_U.if_full_n;
    assign fifo_intf_895.fifo_rd_block = 0;
    assign fifo_intf_895.fifo_wr_block = 0;
    assign fifo_intf_895.finish = finish;
    csv_file_dump fifo_csv_dumper_895;
    csv_file_dump cstatus_csv_dumper_895;
    df_fifo_monitor fifo_monitor_895;
    df_fifo_intf fifo_intf_896(clock,reset);
    assign fifo_intf_896.rd_en = AESL_inst_myproject.layer2_out_895_U.if_read & AESL_inst_myproject.layer2_out_895_U.if_empty_n;
    assign fifo_intf_896.wr_en = AESL_inst_myproject.layer2_out_895_U.if_write & AESL_inst_myproject.layer2_out_895_U.if_full_n;
    assign fifo_intf_896.fifo_rd_block = 0;
    assign fifo_intf_896.fifo_wr_block = 0;
    assign fifo_intf_896.finish = finish;
    csv_file_dump fifo_csv_dumper_896;
    csv_file_dump cstatus_csv_dumper_896;
    df_fifo_monitor fifo_monitor_896;
    df_fifo_intf fifo_intf_897(clock,reset);
    assign fifo_intf_897.rd_en = AESL_inst_myproject.layer2_out_896_U.if_read & AESL_inst_myproject.layer2_out_896_U.if_empty_n;
    assign fifo_intf_897.wr_en = AESL_inst_myproject.layer2_out_896_U.if_write & AESL_inst_myproject.layer2_out_896_U.if_full_n;
    assign fifo_intf_897.fifo_rd_block = 0;
    assign fifo_intf_897.fifo_wr_block = 0;
    assign fifo_intf_897.finish = finish;
    csv_file_dump fifo_csv_dumper_897;
    csv_file_dump cstatus_csv_dumper_897;
    df_fifo_monitor fifo_monitor_897;
    df_fifo_intf fifo_intf_898(clock,reset);
    assign fifo_intf_898.rd_en = AESL_inst_myproject.layer2_out_897_U.if_read & AESL_inst_myproject.layer2_out_897_U.if_empty_n;
    assign fifo_intf_898.wr_en = AESL_inst_myproject.layer2_out_897_U.if_write & AESL_inst_myproject.layer2_out_897_U.if_full_n;
    assign fifo_intf_898.fifo_rd_block = 0;
    assign fifo_intf_898.fifo_wr_block = 0;
    assign fifo_intf_898.finish = finish;
    csv_file_dump fifo_csv_dumper_898;
    csv_file_dump cstatus_csv_dumper_898;
    df_fifo_monitor fifo_monitor_898;
    df_fifo_intf fifo_intf_899(clock,reset);
    assign fifo_intf_899.rd_en = AESL_inst_myproject.layer2_out_898_U.if_read & AESL_inst_myproject.layer2_out_898_U.if_empty_n;
    assign fifo_intf_899.wr_en = AESL_inst_myproject.layer2_out_898_U.if_write & AESL_inst_myproject.layer2_out_898_U.if_full_n;
    assign fifo_intf_899.fifo_rd_block = 0;
    assign fifo_intf_899.fifo_wr_block = 0;
    assign fifo_intf_899.finish = finish;
    csv_file_dump fifo_csv_dumper_899;
    csv_file_dump cstatus_csv_dumper_899;
    df_fifo_monitor fifo_monitor_899;
    df_fifo_intf fifo_intf_900(clock,reset);
    assign fifo_intf_900.rd_en = AESL_inst_myproject.layer2_out_899_U.if_read & AESL_inst_myproject.layer2_out_899_U.if_empty_n;
    assign fifo_intf_900.wr_en = AESL_inst_myproject.layer2_out_899_U.if_write & AESL_inst_myproject.layer2_out_899_U.if_full_n;
    assign fifo_intf_900.fifo_rd_block = 0;
    assign fifo_intf_900.fifo_wr_block = 0;
    assign fifo_intf_900.finish = finish;
    csv_file_dump fifo_csv_dumper_900;
    csv_file_dump cstatus_csv_dumper_900;
    df_fifo_monitor fifo_monitor_900;
    df_fifo_intf fifo_intf_901(clock,reset);
    assign fifo_intf_901.rd_en = AESL_inst_myproject.layer2_out_900_U.if_read & AESL_inst_myproject.layer2_out_900_U.if_empty_n;
    assign fifo_intf_901.wr_en = AESL_inst_myproject.layer2_out_900_U.if_write & AESL_inst_myproject.layer2_out_900_U.if_full_n;
    assign fifo_intf_901.fifo_rd_block = 0;
    assign fifo_intf_901.fifo_wr_block = 0;
    assign fifo_intf_901.finish = finish;
    csv_file_dump fifo_csv_dumper_901;
    csv_file_dump cstatus_csv_dumper_901;
    df_fifo_monitor fifo_monitor_901;
    df_fifo_intf fifo_intf_902(clock,reset);
    assign fifo_intf_902.rd_en = AESL_inst_myproject.layer2_out_901_U.if_read & AESL_inst_myproject.layer2_out_901_U.if_empty_n;
    assign fifo_intf_902.wr_en = AESL_inst_myproject.layer2_out_901_U.if_write & AESL_inst_myproject.layer2_out_901_U.if_full_n;
    assign fifo_intf_902.fifo_rd_block = 0;
    assign fifo_intf_902.fifo_wr_block = 0;
    assign fifo_intf_902.finish = finish;
    csv_file_dump fifo_csv_dumper_902;
    csv_file_dump cstatus_csv_dumper_902;
    df_fifo_monitor fifo_monitor_902;
    df_fifo_intf fifo_intf_903(clock,reset);
    assign fifo_intf_903.rd_en = AESL_inst_myproject.layer2_out_902_U.if_read & AESL_inst_myproject.layer2_out_902_U.if_empty_n;
    assign fifo_intf_903.wr_en = AESL_inst_myproject.layer2_out_902_U.if_write & AESL_inst_myproject.layer2_out_902_U.if_full_n;
    assign fifo_intf_903.fifo_rd_block = 0;
    assign fifo_intf_903.fifo_wr_block = 0;
    assign fifo_intf_903.finish = finish;
    csv_file_dump fifo_csv_dumper_903;
    csv_file_dump cstatus_csv_dumper_903;
    df_fifo_monitor fifo_monitor_903;
    df_fifo_intf fifo_intf_904(clock,reset);
    assign fifo_intf_904.rd_en = AESL_inst_myproject.layer2_out_903_U.if_read & AESL_inst_myproject.layer2_out_903_U.if_empty_n;
    assign fifo_intf_904.wr_en = AESL_inst_myproject.layer2_out_903_U.if_write & AESL_inst_myproject.layer2_out_903_U.if_full_n;
    assign fifo_intf_904.fifo_rd_block = 0;
    assign fifo_intf_904.fifo_wr_block = 0;
    assign fifo_intf_904.finish = finish;
    csv_file_dump fifo_csv_dumper_904;
    csv_file_dump cstatus_csv_dumper_904;
    df_fifo_monitor fifo_monitor_904;
    df_fifo_intf fifo_intf_905(clock,reset);
    assign fifo_intf_905.rd_en = AESL_inst_myproject.layer2_out_904_U.if_read & AESL_inst_myproject.layer2_out_904_U.if_empty_n;
    assign fifo_intf_905.wr_en = AESL_inst_myproject.layer2_out_904_U.if_write & AESL_inst_myproject.layer2_out_904_U.if_full_n;
    assign fifo_intf_905.fifo_rd_block = 0;
    assign fifo_intf_905.fifo_wr_block = 0;
    assign fifo_intf_905.finish = finish;
    csv_file_dump fifo_csv_dumper_905;
    csv_file_dump cstatus_csv_dumper_905;
    df_fifo_monitor fifo_monitor_905;
    df_fifo_intf fifo_intf_906(clock,reset);
    assign fifo_intf_906.rd_en = AESL_inst_myproject.layer2_out_905_U.if_read & AESL_inst_myproject.layer2_out_905_U.if_empty_n;
    assign fifo_intf_906.wr_en = AESL_inst_myproject.layer2_out_905_U.if_write & AESL_inst_myproject.layer2_out_905_U.if_full_n;
    assign fifo_intf_906.fifo_rd_block = 0;
    assign fifo_intf_906.fifo_wr_block = 0;
    assign fifo_intf_906.finish = finish;
    csv_file_dump fifo_csv_dumper_906;
    csv_file_dump cstatus_csv_dumper_906;
    df_fifo_monitor fifo_monitor_906;
    df_fifo_intf fifo_intf_907(clock,reset);
    assign fifo_intf_907.rd_en = AESL_inst_myproject.layer2_out_906_U.if_read & AESL_inst_myproject.layer2_out_906_U.if_empty_n;
    assign fifo_intf_907.wr_en = AESL_inst_myproject.layer2_out_906_U.if_write & AESL_inst_myproject.layer2_out_906_U.if_full_n;
    assign fifo_intf_907.fifo_rd_block = 0;
    assign fifo_intf_907.fifo_wr_block = 0;
    assign fifo_intf_907.finish = finish;
    csv_file_dump fifo_csv_dumper_907;
    csv_file_dump cstatus_csv_dumper_907;
    df_fifo_monitor fifo_monitor_907;
    df_fifo_intf fifo_intf_908(clock,reset);
    assign fifo_intf_908.rd_en = AESL_inst_myproject.layer2_out_907_U.if_read & AESL_inst_myproject.layer2_out_907_U.if_empty_n;
    assign fifo_intf_908.wr_en = AESL_inst_myproject.layer2_out_907_U.if_write & AESL_inst_myproject.layer2_out_907_U.if_full_n;
    assign fifo_intf_908.fifo_rd_block = 0;
    assign fifo_intf_908.fifo_wr_block = 0;
    assign fifo_intf_908.finish = finish;
    csv_file_dump fifo_csv_dumper_908;
    csv_file_dump cstatus_csv_dumper_908;
    df_fifo_monitor fifo_monitor_908;
    df_fifo_intf fifo_intf_909(clock,reset);
    assign fifo_intf_909.rd_en = AESL_inst_myproject.layer2_out_908_U.if_read & AESL_inst_myproject.layer2_out_908_U.if_empty_n;
    assign fifo_intf_909.wr_en = AESL_inst_myproject.layer2_out_908_U.if_write & AESL_inst_myproject.layer2_out_908_U.if_full_n;
    assign fifo_intf_909.fifo_rd_block = 0;
    assign fifo_intf_909.fifo_wr_block = 0;
    assign fifo_intf_909.finish = finish;
    csv_file_dump fifo_csv_dumper_909;
    csv_file_dump cstatus_csv_dumper_909;
    df_fifo_monitor fifo_monitor_909;
    df_fifo_intf fifo_intf_910(clock,reset);
    assign fifo_intf_910.rd_en = AESL_inst_myproject.layer2_out_909_U.if_read & AESL_inst_myproject.layer2_out_909_U.if_empty_n;
    assign fifo_intf_910.wr_en = AESL_inst_myproject.layer2_out_909_U.if_write & AESL_inst_myproject.layer2_out_909_U.if_full_n;
    assign fifo_intf_910.fifo_rd_block = 0;
    assign fifo_intf_910.fifo_wr_block = 0;
    assign fifo_intf_910.finish = finish;
    csv_file_dump fifo_csv_dumper_910;
    csv_file_dump cstatus_csv_dumper_910;
    df_fifo_monitor fifo_monitor_910;
    df_fifo_intf fifo_intf_911(clock,reset);
    assign fifo_intf_911.rd_en = AESL_inst_myproject.layer2_out_910_U.if_read & AESL_inst_myproject.layer2_out_910_U.if_empty_n;
    assign fifo_intf_911.wr_en = AESL_inst_myproject.layer2_out_910_U.if_write & AESL_inst_myproject.layer2_out_910_U.if_full_n;
    assign fifo_intf_911.fifo_rd_block = 0;
    assign fifo_intf_911.fifo_wr_block = 0;
    assign fifo_intf_911.finish = finish;
    csv_file_dump fifo_csv_dumper_911;
    csv_file_dump cstatus_csv_dumper_911;
    df_fifo_monitor fifo_monitor_911;
    df_fifo_intf fifo_intf_912(clock,reset);
    assign fifo_intf_912.rd_en = AESL_inst_myproject.layer2_out_911_U.if_read & AESL_inst_myproject.layer2_out_911_U.if_empty_n;
    assign fifo_intf_912.wr_en = AESL_inst_myproject.layer2_out_911_U.if_write & AESL_inst_myproject.layer2_out_911_U.if_full_n;
    assign fifo_intf_912.fifo_rd_block = 0;
    assign fifo_intf_912.fifo_wr_block = 0;
    assign fifo_intf_912.finish = finish;
    csv_file_dump fifo_csv_dumper_912;
    csv_file_dump cstatus_csv_dumper_912;
    df_fifo_monitor fifo_monitor_912;
    df_fifo_intf fifo_intf_913(clock,reset);
    assign fifo_intf_913.rd_en = AESL_inst_myproject.layer2_out_912_U.if_read & AESL_inst_myproject.layer2_out_912_U.if_empty_n;
    assign fifo_intf_913.wr_en = AESL_inst_myproject.layer2_out_912_U.if_write & AESL_inst_myproject.layer2_out_912_U.if_full_n;
    assign fifo_intf_913.fifo_rd_block = 0;
    assign fifo_intf_913.fifo_wr_block = 0;
    assign fifo_intf_913.finish = finish;
    csv_file_dump fifo_csv_dumper_913;
    csv_file_dump cstatus_csv_dumper_913;
    df_fifo_monitor fifo_monitor_913;
    df_fifo_intf fifo_intf_914(clock,reset);
    assign fifo_intf_914.rd_en = AESL_inst_myproject.layer2_out_913_U.if_read & AESL_inst_myproject.layer2_out_913_U.if_empty_n;
    assign fifo_intf_914.wr_en = AESL_inst_myproject.layer2_out_913_U.if_write & AESL_inst_myproject.layer2_out_913_U.if_full_n;
    assign fifo_intf_914.fifo_rd_block = 0;
    assign fifo_intf_914.fifo_wr_block = 0;
    assign fifo_intf_914.finish = finish;
    csv_file_dump fifo_csv_dumper_914;
    csv_file_dump cstatus_csv_dumper_914;
    df_fifo_monitor fifo_monitor_914;
    df_fifo_intf fifo_intf_915(clock,reset);
    assign fifo_intf_915.rd_en = AESL_inst_myproject.layer2_out_914_U.if_read & AESL_inst_myproject.layer2_out_914_U.if_empty_n;
    assign fifo_intf_915.wr_en = AESL_inst_myproject.layer2_out_914_U.if_write & AESL_inst_myproject.layer2_out_914_U.if_full_n;
    assign fifo_intf_915.fifo_rd_block = 0;
    assign fifo_intf_915.fifo_wr_block = 0;
    assign fifo_intf_915.finish = finish;
    csv_file_dump fifo_csv_dumper_915;
    csv_file_dump cstatus_csv_dumper_915;
    df_fifo_monitor fifo_monitor_915;
    df_fifo_intf fifo_intf_916(clock,reset);
    assign fifo_intf_916.rd_en = AESL_inst_myproject.layer2_out_915_U.if_read & AESL_inst_myproject.layer2_out_915_U.if_empty_n;
    assign fifo_intf_916.wr_en = AESL_inst_myproject.layer2_out_915_U.if_write & AESL_inst_myproject.layer2_out_915_U.if_full_n;
    assign fifo_intf_916.fifo_rd_block = 0;
    assign fifo_intf_916.fifo_wr_block = 0;
    assign fifo_intf_916.finish = finish;
    csv_file_dump fifo_csv_dumper_916;
    csv_file_dump cstatus_csv_dumper_916;
    df_fifo_monitor fifo_monitor_916;
    df_fifo_intf fifo_intf_917(clock,reset);
    assign fifo_intf_917.rd_en = AESL_inst_myproject.layer2_out_916_U.if_read & AESL_inst_myproject.layer2_out_916_U.if_empty_n;
    assign fifo_intf_917.wr_en = AESL_inst_myproject.layer2_out_916_U.if_write & AESL_inst_myproject.layer2_out_916_U.if_full_n;
    assign fifo_intf_917.fifo_rd_block = 0;
    assign fifo_intf_917.fifo_wr_block = 0;
    assign fifo_intf_917.finish = finish;
    csv_file_dump fifo_csv_dumper_917;
    csv_file_dump cstatus_csv_dumper_917;
    df_fifo_monitor fifo_monitor_917;
    df_fifo_intf fifo_intf_918(clock,reset);
    assign fifo_intf_918.rd_en = AESL_inst_myproject.layer2_out_917_U.if_read & AESL_inst_myproject.layer2_out_917_U.if_empty_n;
    assign fifo_intf_918.wr_en = AESL_inst_myproject.layer2_out_917_U.if_write & AESL_inst_myproject.layer2_out_917_U.if_full_n;
    assign fifo_intf_918.fifo_rd_block = 0;
    assign fifo_intf_918.fifo_wr_block = 0;
    assign fifo_intf_918.finish = finish;
    csv_file_dump fifo_csv_dumper_918;
    csv_file_dump cstatus_csv_dumper_918;
    df_fifo_monitor fifo_monitor_918;
    df_fifo_intf fifo_intf_919(clock,reset);
    assign fifo_intf_919.rd_en = AESL_inst_myproject.layer2_out_918_U.if_read & AESL_inst_myproject.layer2_out_918_U.if_empty_n;
    assign fifo_intf_919.wr_en = AESL_inst_myproject.layer2_out_918_U.if_write & AESL_inst_myproject.layer2_out_918_U.if_full_n;
    assign fifo_intf_919.fifo_rd_block = 0;
    assign fifo_intf_919.fifo_wr_block = 0;
    assign fifo_intf_919.finish = finish;
    csv_file_dump fifo_csv_dumper_919;
    csv_file_dump cstatus_csv_dumper_919;
    df_fifo_monitor fifo_monitor_919;
    df_fifo_intf fifo_intf_920(clock,reset);
    assign fifo_intf_920.rd_en = AESL_inst_myproject.layer2_out_919_U.if_read & AESL_inst_myproject.layer2_out_919_U.if_empty_n;
    assign fifo_intf_920.wr_en = AESL_inst_myproject.layer2_out_919_U.if_write & AESL_inst_myproject.layer2_out_919_U.if_full_n;
    assign fifo_intf_920.fifo_rd_block = 0;
    assign fifo_intf_920.fifo_wr_block = 0;
    assign fifo_intf_920.finish = finish;
    csv_file_dump fifo_csv_dumper_920;
    csv_file_dump cstatus_csv_dumper_920;
    df_fifo_monitor fifo_monitor_920;
    df_fifo_intf fifo_intf_921(clock,reset);
    assign fifo_intf_921.rd_en = AESL_inst_myproject.layer2_out_920_U.if_read & AESL_inst_myproject.layer2_out_920_U.if_empty_n;
    assign fifo_intf_921.wr_en = AESL_inst_myproject.layer2_out_920_U.if_write & AESL_inst_myproject.layer2_out_920_U.if_full_n;
    assign fifo_intf_921.fifo_rd_block = 0;
    assign fifo_intf_921.fifo_wr_block = 0;
    assign fifo_intf_921.finish = finish;
    csv_file_dump fifo_csv_dumper_921;
    csv_file_dump cstatus_csv_dumper_921;
    df_fifo_monitor fifo_monitor_921;
    df_fifo_intf fifo_intf_922(clock,reset);
    assign fifo_intf_922.rd_en = AESL_inst_myproject.layer2_out_921_U.if_read & AESL_inst_myproject.layer2_out_921_U.if_empty_n;
    assign fifo_intf_922.wr_en = AESL_inst_myproject.layer2_out_921_U.if_write & AESL_inst_myproject.layer2_out_921_U.if_full_n;
    assign fifo_intf_922.fifo_rd_block = 0;
    assign fifo_intf_922.fifo_wr_block = 0;
    assign fifo_intf_922.finish = finish;
    csv_file_dump fifo_csv_dumper_922;
    csv_file_dump cstatus_csv_dumper_922;
    df_fifo_monitor fifo_monitor_922;
    df_fifo_intf fifo_intf_923(clock,reset);
    assign fifo_intf_923.rd_en = AESL_inst_myproject.layer2_out_922_U.if_read & AESL_inst_myproject.layer2_out_922_U.if_empty_n;
    assign fifo_intf_923.wr_en = AESL_inst_myproject.layer2_out_922_U.if_write & AESL_inst_myproject.layer2_out_922_U.if_full_n;
    assign fifo_intf_923.fifo_rd_block = 0;
    assign fifo_intf_923.fifo_wr_block = 0;
    assign fifo_intf_923.finish = finish;
    csv_file_dump fifo_csv_dumper_923;
    csv_file_dump cstatus_csv_dumper_923;
    df_fifo_monitor fifo_monitor_923;
    df_fifo_intf fifo_intf_924(clock,reset);
    assign fifo_intf_924.rd_en = AESL_inst_myproject.layer2_out_923_U.if_read & AESL_inst_myproject.layer2_out_923_U.if_empty_n;
    assign fifo_intf_924.wr_en = AESL_inst_myproject.layer2_out_923_U.if_write & AESL_inst_myproject.layer2_out_923_U.if_full_n;
    assign fifo_intf_924.fifo_rd_block = 0;
    assign fifo_intf_924.fifo_wr_block = 0;
    assign fifo_intf_924.finish = finish;
    csv_file_dump fifo_csv_dumper_924;
    csv_file_dump cstatus_csv_dumper_924;
    df_fifo_monitor fifo_monitor_924;
    df_fifo_intf fifo_intf_925(clock,reset);
    assign fifo_intf_925.rd_en = AESL_inst_myproject.layer2_out_924_U.if_read & AESL_inst_myproject.layer2_out_924_U.if_empty_n;
    assign fifo_intf_925.wr_en = AESL_inst_myproject.layer2_out_924_U.if_write & AESL_inst_myproject.layer2_out_924_U.if_full_n;
    assign fifo_intf_925.fifo_rd_block = 0;
    assign fifo_intf_925.fifo_wr_block = 0;
    assign fifo_intf_925.finish = finish;
    csv_file_dump fifo_csv_dumper_925;
    csv_file_dump cstatus_csv_dumper_925;
    df_fifo_monitor fifo_monitor_925;
    df_fifo_intf fifo_intf_926(clock,reset);
    assign fifo_intf_926.rd_en = AESL_inst_myproject.layer2_out_925_U.if_read & AESL_inst_myproject.layer2_out_925_U.if_empty_n;
    assign fifo_intf_926.wr_en = AESL_inst_myproject.layer2_out_925_U.if_write & AESL_inst_myproject.layer2_out_925_U.if_full_n;
    assign fifo_intf_926.fifo_rd_block = 0;
    assign fifo_intf_926.fifo_wr_block = 0;
    assign fifo_intf_926.finish = finish;
    csv_file_dump fifo_csv_dumper_926;
    csv_file_dump cstatus_csv_dumper_926;
    df_fifo_monitor fifo_monitor_926;
    df_fifo_intf fifo_intf_927(clock,reset);
    assign fifo_intf_927.rd_en = AESL_inst_myproject.layer2_out_926_U.if_read & AESL_inst_myproject.layer2_out_926_U.if_empty_n;
    assign fifo_intf_927.wr_en = AESL_inst_myproject.layer2_out_926_U.if_write & AESL_inst_myproject.layer2_out_926_U.if_full_n;
    assign fifo_intf_927.fifo_rd_block = 0;
    assign fifo_intf_927.fifo_wr_block = 0;
    assign fifo_intf_927.finish = finish;
    csv_file_dump fifo_csv_dumper_927;
    csv_file_dump cstatus_csv_dumper_927;
    df_fifo_monitor fifo_monitor_927;
    df_fifo_intf fifo_intf_928(clock,reset);
    assign fifo_intf_928.rd_en = AESL_inst_myproject.layer2_out_927_U.if_read & AESL_inst_myproject.layer2_out_927_U.if_empty_n;
    assign fifo_intf_928.wr_en = AESL_inst_myproject.layer2_out_927_U.if_write & AESL_inst_myproject.layer2_out_927_U.if_full_n;
    assign fifo_intf_928.fifo_rd_block = 0;
    assign fifo_intf_928.fifo_wr_block = 0;
    assign fifo_intf_928.finish = finish;
    csv_file_dump fifo_csv_dumper_928;
    csv_file_dump cstatus_csv_dumper_928;
    df_fifo_monitor fifo_monitor_928;
    df_fifo_intf fifo_intf_929(clock,reset);
    assign fifo_intf_929.rd_en = AESL_inst_myproject.layer2_out_928_U.if_read & AESL_inst_myproject.layer2_out_928_U.if_empty_n;
    assign fifo_intf_929.wr_en = AESL_inst_myproject.layer2_out_928_U.if_write & AESL_inst_myproject.layer2_out_928_U.if_full_n;
    assign fifo_intf_929.fifo_rd_block = 0;
    assign fifo_intf_929.fifo_wr_block = 0;
    assign fifo_intf_929.finish = finish;
    csv_file_dump fifo_csv_dumper_929;
    csv_file_dump cstatus_csv_dumper_929;
    df_fifo_monitor fifo_monitor_929;
    df_fifo_intf fifo_intf_930(clock,reset);
    assign fifo_intf_930.rd_en = AESL_inst_myproject.layer2_out_929_U.if_read & AESL_inst_myproject.layer2_out_929_U.if_empty_n;
    assign fifo_intf_930.wr_en = AESL_inst_myproject.layer2_out_929_U.if_write & AESL_inst_myproject.layer2_out_929_U.if_full_n;
    assign fifo_intf_930.fifo_rd_block = 0;
    assign fifo_intf_930.fifo_wr_block = 0;
    assign fifo_intf_930.finish = finish;
    csv_file_dump fifo_csv_dumper_930;
    csv_file_dump cstatus_csv_dumper_930;
    df_fifo_monitor fifo_monitor_930;
    df_fifo_intf fifo_intf_931(clock,reset);
    assign fifo_intf_931.rd_en = AESL_inst_myproject.layer2_out_930_U.if_read & AESL_inst_myproject.layer2_out_930_U.if_empty_n;
    assign fifo_intf_931.wr_en = AESL_inst_myproject.layer2_out_930_U.if_write & AESL_inst_myproject.layer2_out_930_U.if_full_n;
    assign fifo_intf_931.fifo_rd_block = 0;
    assign fifo_intf_931.fifo_wr_block = 0;
    assign fifo_intf_931.finish = finish;
    csv_file_dump fifo_csv_dumper_931;
    csv_file_dump cstatus_csv_dumper_931;
    df_fifo_monitor fifo_monitor_931;
    df_fifo_intf fifo_intf_932(clock,reset);
    assign fifo_intf_932.rd_en = AESL_inst_myproject.layer2_out_931_U.if_read & AESL_inst_myproject.layer2_out_931_U.if_empty_n;
    assign fifo_intf_932.wr_en = AESL_inst_myproject.layer2_out_931_U.if_write & AESL_inst_myproject.layer2_out_931_U.if_full_n;
    assign fifo_intf_932.fifo_rd_block = 0;
    assign fifo_intf_932.fifo_wr_block = 0;
    assign fifo_intf_932.finish = finish;
    csv_file_dump fifo_csv_dumper_932;
    csv_file_dump cstatus_csv_dumper_932;
    df_fifo_monitor fifo_monitor_932;
    df_fifo_intf fifo_intf_933(clock,reset);
    assign fifo_intf_933.rd_en = AESL_inst_myproject.layer2_out_932_U.if_read & AESL_inst_myproject.layer2_out_932_U.if_empty_n;
    assign fifo_intf_933.wr_en = AESL_inst_myproject.layer2_out_932_U.if_write & AESL_inst_myproject.layer2_out_932_U.if_full_n;
    assign fifo_intf_933.fifo_rd_block = 0;
    assign fifo_intf_933.fifo_wr_block = 0;
    assign fifo_intf_933.finish = finish;
    csv_file_dump fifo_csv_dumper_933;
    csv_file_dump cstatus_csv_dumper_933;
    df_fifo_monitor fifo_monitor_933;
    df_fifo_intf fifo_intf_934(clock,reset);
    assign fifo_intf_934.rd_en = AESL_inst_myproject.layer2_out_933_U.if_read & AESL_inst_myproject.layer2_out_933_U.if_empty_n;
    assign fifo_intf_934.wr_en = AESL_inst_myproject.layer2_out_933_U.if_write & AESL_inst_myproject.layer2_out_933_U.if_full_n;
    assign fifo_intf_934.fifo_rd_block = 0;
    assign fifo_intf_934.fifo_wr_block = 0;
    assign fifo_intf_934.finish = finish;
    csv_file_dump fifo_csv_dumper_934;
    csv_file_dump cstatus_csv_dumper_934;
    df_fifo_monitor fifo_monitor_934;
    df_fifo_intf fifo_intf_935(clock,reset);
    assign fifo_intf_935.rd_en = AESL_inst_myproject.layer2_out_934_U.if_read & AESL_inst_myproject.layer2_out_934_U.if_empty_n;
    assign fifo_intf_935.wr_en = AESL_inst_myproject.layer2_out_934_U.if_write & AESL_inst_myproject.layer2_out_934_U.if_full_n;
    assign fifo_intf_935.fifo_rd_block = 0;
    assign fifo_intf_935.fifo_wr_block = 0;
    assign fifo_intf_935.finish = finish;
    csv_file_dump fifo_csv_dumper_935;
    csv_file_dump cstatus_csv_dumper_935;
    df_fifo_monitor fifo_monitor_935;
    df_fifo_intf fifo_intf_936(clock,reset);
    assign fifo_intf_936.rd_en = AESL_inst_myproject.layer2_out_935_U.if_read & AESL_inst_myproject.layer2_out_935_U.if_empty_n;
    assign fifo_intf_936.wr_en = AESL_inst_myproject.layer2_out_935_U.if_write & AESL_inst_myproject.layer2_out_935_U.if_full_n;
    assign fifo_intf_936.fifo_rd_block = 0;
    assign fifo_intf_936.fifo_wr_block = 0;
    assign fifo_intf_936.finish = finish;
    csv_file_dump fifo_csv_dumper_936;
    csv_file_dump cstatus_csv_dumper_936;
    df_fifo_monitor fifo_monitor_936;
    df_fifo_intf fifo_intf_937(clock,reset);
    assign fifo_intf_937.rd_en = AESL_inst_myproject.layer2_out_936_U.if_read & AESL_inst_myproject.layer2_out_936_U.if_empty_n;
    assign fifo_intf_937.wr_en = AESL_inst_myproject.layer2_out_936_U.if_write & AESL_inst_myproject.layer2_out_936_U.if_full_n;
    assign fifo_intf_937.fifo_rd_block = 0;
    assign fifo_intf_937.fifo_wr_block = 0;
    assign fifo_intf_937.finish = finish;
    csv_file_dump fifo_csv_dumper_937;
    csv_file_dump cstatus_csv_dumper_937;
    df_fifo_monitor fifo_monitor_937;
    df_fifo_intf fifo_intf_938(clock,reset);
    assign fifo_intf_938.rd_en = AESL_inst_myproject.layer2_out_937_U.if_read & AESL_inst_myproject.layer2_out_937_U.if_empty_n;
    assign fifo_intf_938.wr_en = AESL_inst_myproject.layer2_out_937_U.if_write & AESL_inst_myproject.layer2_out_937_U.if_full_n;
    assign fifo_intf_938.fifo_rd_block = 0;
    assign fifo_intf_938.fifo_wr_block = 0;
    assign fifo_intf_938.finish = finish;
    csv_file_dump fifo_csv_dumper_938;
    csv_file_dump cstatus_csv_dumper_938;
    df_fifo_monitor fifo_monitor_938;
    df_fifo_intf fifo_intf_939(clock,reset);
    assign fifo_intf_939.rd_en = AESL_inst_myproject.layer2_out_938_U.if_read & AESL_inst_myproject.layer2_out_938_U.if_empty_n;
    assign fifo_intf_939.wr_en = AESL_inst_myproject.layer2_out_938_U.if_write & AESL_inst_myproject.layer2_out_938_U.if_full_n;
    assign fifo_intf_939.fifo_rd_block = 0;
    assign fifo_intf_939.fifo_wr_block = 0;
    assign fifo_intf_939.finish = finish;
    csv_file_dump fifo_csv_dumper_939;
    csv_file_dump cstatus_csv_dumper_939;
    df_fifo_monitor fifo_monitor_939;
    df_fifo_intf fifo_intf_940(clock,reset);
    assign fifo_intf_940.rd_en = AESL_inst_myproject.layer2_out_939_U.if_read & AESL_inst_myproject.layer2_out_939_U.if_empty_n;
    assign fifo_intf_940.wr_en = AESL_inst_myproject.layer2_out_939_U.if_write & AESL_inst_myproject.layer2_out_939_U.if_full_n;
    assign fifo_intf_940.fifo_rd_block = 0;
    assign fifo_intf_940.fifo_wr_block = 0;
    assign fifo_intf_940.finish = finish;
    csv_file_dump fifo_csv_dumper_940;
    csv_file_dump cstatus_csv_dumper_940;
    df_fifo_monitor fifo_monitor_940;
    df_fifo_intf fifo_intf_941(clock,reset);
    assign fifo_intf_941.rd_en = AESL_inst_myproject.layer2_out_940_U.if_read & AESL_inst_myproject.layer2_out_940_U.if_empty_n;
    assign fifo_intf_941.wr_en = AESL_inst_myproject.layer2_out_940_U.if_write & AESL_inst_myproject.layer2_out_940_U.if_full_n;
    assign fifo_intf_941.fifo_rd_block = 0;
    assign fifo_intf_941.fifo_wr_block = 0;
    assign fifo_intf_941.finish = finish;
    csv_file_dump fifo_csv_dumper_941;
    csv_file_dump cstatus_csv_dumper_941;
    df_fifo_monitor fifo_monitor_941;
    df_fifo_intf fifo_intf_942(clock,reset);
    assign fifo_intf_942.rd_en = AESL_inst_myproject.layer2_out_941_U.if_read & AESL_inst_myproject.layer2_out_941_U.if_empty_n;
    assign fifo_intf_942.wr_en = AESL_inst_myproject.layer2_out_941_U.if_write & AESL_inst_myproject.layer2_out_941_U.if_full_n;
    assign fifo_intf_942.fifo_rd_block = 0;
    assign fifo_intf_942.fifo_wr_block = 0;
    assign fifo_intf_942.finish = finish;
    csv_file_dump fifo_csv_dumper_942;
    csv_file_dump cstatus_csv_dumper_942;
    df_fifo_monitor fifo_monitor_942;
    df_fifo_intf fifo_intf_943(clock,reset);
    assign fifo_intf_943.rd_en = AESL_inst_myproject.layer2_out_942_U.if_read & AESL_inst_myproject.layer2_out_942_U.if_empty_n;
    assign fifo_intf_943.wr_en = AESL_inst_myproject.layer2_out_942_U.if_write & AESL_inst_myproject.layer2_out_942_U.if_full_n;
    assign fifo_intf_943.fifo_rd_block = 0;
    assign fifo_intf_943.fifo_wr_block = 0;
    assign fifo_intf_943.finish = finish;
    csv_file_dump fifo_csv_dumper_943;
    csv_file_dump cstatus_csv_dumper_943;
    df_fifo_monitor fifo_monitor_943;
    df_fifo_intf fifo_intf_944(clock,reset);
    assign fifo_intf_944.rd_en = AESL_inst_myproject.layer2_out_943_U.if_read & AESL_inst_myproject.layer2_out_943_U.if_empty_n;
    assign fifo_intf_944.wr_en = AESL_inst_myproject.layer2_out_943_U.if_write & AESL_inst_myproject.layer2_out_943_U.if_full_n;
    assign fifo_intf_944.fifo_rd_block = 0;
    assign fifo_intf_944.fifo_wr_block = 0;
    assign fifo_intf_944.finish = finish;
    csv_file_dump fifo_csv_dumper_944;
    csv_file_dump cstatus_csv_dumper_944;
    df_fifo_monitor fifo_monitor_944;
    df_fifo_intf fifo_intf_945(clock,reset);
    assign fifo_intf_945.rd_en = AESL_inst_myproject.layer2_out_944_U.if_read & AESL_inst_myproject.layer2_out_944_U.if_empty_n;
    assign fifo_intf_945.wr_en = AESL_inst_myproject.layer2_out_944_U.if_write & AESL_inst_myproject.layer2_out_944_U.if_full_n;
    assign fifo_intf_945.fifo_rd_block = 0;
    assign fifo_intf_945.fifo_wr_block = 0;
    assign fifo_intf_945.finish = finish;
    csv_file_dump fifo_csv_dumper_945;
    csv_file_dump cstatus_csv_dumper_945;
    df_fifo_monitor fifo_monitor_945;
    df_fifo_intf fifo_intf_946(clock,reset);
    assign fifo_intf_946.rd_en = AESL_inst_myproject.layer2_out_945_U.if_read & AESL_inst_myproject.layer2_out_945_U.if_empty_n;
    assign fifo_intf_946.wr_en = AESL_inst_myproject.layer2_out_945_U.if_write & AESL_inst_myproject.layer2_out_945_U.if_full_n;
    assign fifo_intf_946.fifo_rd_block = 0;
    assign fifo_intf_946.fifo_wr_block = 0;
    assign fifo_intf_946.finish = finish;
    csv_file_dump fifo_csv_dumper_946;
    csv_file_dump cstatus_csv_dumper_946;
    df_fifo_monitor fifo_monitor_946;
    df_fifo_intf fifo_intf_947(clock,reset);
    assign fifo_intf_947.rd_en = AESL_inst_myproject.layer2_out_946_U.if_read & AESL_inst_myproject.layer2_out_946_U.if_empty_n;
    assign fifo_intf_947.wr_en = AESL_inst_myproject.layer2_out_946_U.if_write & AESL_inst_myproject.layer2_out_946_U.if_full_n;
    assign fifo_intf_947.fifo_rd_block = 0;
    assign fifo_intf_947.fifo_wr_block = 0;
    assign fifo_intf_947.finish = finish;
    csv_file_dump fifo_csv_dumper_947;
    csv_file_dump cstatus_csv_dumper_947;
    df_fifo_monitor fifo_monitor_947;
    df_fifo_intf fifo_intf_948(clock,reset);
    assign fifo_intf_948.rd_en = AESL_inst_myproject.layer2_out_947_U.if_read & AESL_inst_myproject.layer2_out_947_U.if_empty_n;
    assign fifo_intf_948.wr_en = AESL_inst_myproject.layer2_out_947_U.if_write & AESL_inst_myproject.layer2_out_947_U.if_full_n;
    assign fifo_intf_948.fifo_rd_block = 0;
    assign fifo_intf_948.fifo_wr_block = 0;
    assign fifo_intf_948.finish = finish;
    csv_file_dump fifo_csv_dumper_948;
    csv_file_dump cstatus_csv_dumper_948;
    df_fifo_monitor fifo_monitor_948;
    df_fifo_intf fifo_intf_949(clock,reset);
    assign fifo_intf_949.rd_en = AESL_inst_myproject.layer2_out_948_U.if_read & AESL_inst_myproject.layer2_out_948_U.if_empty_n;
    assign fifo_intf_949.wr_en = AESL_inst_myproject.layer2_out_948_U.if_write & AESL_inst_myproject.layer2_out_948_U.if_full_n;
    assign fifo_intf_949.fifo_rd_block = 0;
    assign fifo_intf_949.fifo_wr_block = 0;
    assign fifo_intf_949.finish = finish;
    csv_file_dump fifo_csv_dumper_949;
    csv_file_dump cstatus_csv_dumper_949;
    df_fifo_monitor fifo_monitor_949;
    df_fifo_intf fifo_intf_950(clock,reset);
    assign fifo_intf_950.rd_en = AESL_inst_myproject.layer2_out_949_U.if_read & AESL_inst_myproject.layer2_out_949_U.if_empty_n;
    assign fifo_intf_950.wr_en = AESL_inst_myproject.layer2_out_949_U.if_write & AESL_inst_myproject.layer2_out_949_U.if_full_n;
    assign fifo_intf_950.fifo_rd_block = 0;
    assign fifo_intf_950.fifo_wr_block = 0;
    assign fifo_intf_950.finish = finish;
    csv_file_dump fifo_csv_dumper_950;
    csv_file_dump cstatus_csv_dumper_950;
    df_fifo_monitor fifo_monitor_950;
    df_fifo_intf fifo_intf_951(clock,reset);
    assign fifo_intf_951.rd_en = AESL_inst_myproject.layer2_out_950_U.if_read & AESL_inst_myproject.layer2_out_950_U.if_empty_n;
    assign fifo_intf_951.wr_en = AESL_inst_myproject.layer2_out_950_U.if_write & AESL_inst_myproject.layer2_out_950_U.if_full_n;
    assign fifo_intf_951.fifo_rd_block = 0;
    assign fifo_intf_951.fifo_wr_block = 0;
    assign fifo_intf_951.finish = finish;
    csv_file_dump fifo_csv_dumper_951;
    csv_file_dump cstatus_csv_dumper_951;
    df_fifo_monitor fifo_monitor_951;
    df_fifo_intf fifo_intf_952(clock,reset);
    assign fifo_intf_952.rd_en = AESL_inst_myproject.layer2_out_951_U.if_read & AESL_inst_myproject.layer2_out_951_U.if_empty_n;
    assign fifo_intf_952.wr_en = AESL_inst_myproject.layer2_out_951_U.if_write & AESL_inst_myproject.layer2_out_951_U.if_full_n;
    assign fifo_intf_952.fifo_rd_block = 0;
    assign fifo_intf_952.fifo_wr_block = 0;
    assign fifo_intf_952.finish = finish;
    csv_file_dump fifo_csv_dumper_952;
    csv_file_dump cstatus_csv_dumper_952;
    df_fifo_monitor fifo_monitor_952;
    df_fifo_intf fifo_intf_953(clock,reset);
    assign fifo_intf_953.rd_en = AESL_inst_myproject.layer2_out_952_U.if_read & AESL_inst_myproject.layer2_out_952_U.if_empty_n;
    assign fifo_intf_953.wr_en = AESL_inst_myproject.layer2_out_952_U.if_write & AESL_inst_myproject.layer2_out_952_U.if_full_n;
    assign fifo_intf_953.fifo_rd_block = 0;
    assign fifo_intf_953.fifo_wr_block = 0;
    assign fifo_intf_953.finish = finish;
    csv_file_dump fifo_csv_dumper_953;
    csv_file_dump cstatus_csv_dumper_953;
    df_fifo_monitor fifo_monitor_953;
    df_fifo_intf fifo_intf_954(clock,reset);
    assign fifo_intf_954.rd_en = AESL_inst_myproject.layer2_out_953_U.if_read & AESL_inst_myproject.layer2_out_953_U.if_empty_n;
    assign fifo_intf_954.wr_en = AESL_inst_myproject.layer2_out_953_U.if_write & AESL_inst_myproject.layer2_out_953_U.if_full_n;
    assign fifo_intf_954.fifo_rd_block = 0;
    assign fifo_intf_954.fifo_wr_block = 0;
    assign fifo_intf_954.finish = finish;
    csv_file_dump fifo_csv_dumper_954;
    csv_file_dump cstatus_csv_dumper_954;
    df_fifo_monitor fifo_monitor_954;
    df_fifo_intf fifo_intf_955(clock,reset);
    assign fifo_intf_955.rd_en = AESL_inst_myproject.layer2_out_954_U.if_read & AESL_inst_myproject.layer2_out_954_U.if_empty_n;
    assign fifo_intf_955.wr_en = AESL_inst_myproject.layer2_out_954_U.if_write & AESL_inst_myproject.layer2_out_954_U.if_full_n;
    assign fifo_intf_955.fifo_rd_block = 0;
    assign fifo_intf_955.fifo_wr_block = 0;
    assign fifo_intf_955.finish = finish;
    csv_file_dump fifo_csv_dumper_955;
    csv_file_dump cstatus_csv_dumper_955;
    df_fifo_monitor fifo_monitor_955;
    df_fifo_intf fifo_intf_956(clock,reset);
    assign fifo_intf_956.rd_en = AESL_inst_myproject.layer2_out_955_U.if_read & AESL_inst_myproject.layer2_out_955_U.if_empty_n;
    assign fifo_intf_956.wr_en = AESL_inst_myproject.layer2_out_955_U.if_write & AESL_inst_myproject.layer2_out_955_U.if_full_n;
    assign fifo_intf_956.fifo_rd_block = 0;
    assign fifo_intf_956.fifo_wr_block = 0;
    assign fifo_intf_956.finish = finish;
    csv_file_dump fifo_csv_dumper_956;
    csv_file_dump cstatus_csv_dumper_956;
    df_fifo_monitor fifo_monitor_956;
    df_fifo_intf fifo_intf_957(clock,reset);
    assign fifo_intf_957.rd_en = AESL_inst_myproject.layer2_out_956_U.if_read & AESL_inst_myproject.layer2_out_956_U.if_empty_n;
    assign fifo_intf_957.wr_en = AESL_inst_myproject.layer2_out_956_U.if_write & AESL_inst_myproject.layer2_out_956_U.if_full_n;
    assign fifo_intf_957.fifo_rd_block = 0;
    assign fifo_intf_957.fifo_wr_block = 0;
    assign fifo_intf_957.finish = finish;
    csv_file_dump fifo_csv_dumper_957;
    csv_file_dump cstatus_csv_dumper_957;
    df_fifo_monitor fifo_monitor_957;
    df_fifo_intf fifo_intf_958(clock,reset);
    assign fifo_intf_958.rd_en = AESL_inst_myproject.layer2_out_957_U.if_read & AESL_inst_myproject.layer2_out_957_U.if_empty_n;
    assign fifo_intf_958.wr_en = AESL_inst_myproject.layer2_out_957_U.if_write & AESL_inst_myproject.layer2_out_957_U.if_full_n;
    assign fifo_intf_958.fifo_rd_block = 0;
    assign fifo_intf_958.fifo_wr_block = 0;
    assign fifo_intf_958.finish = finish;
    csv_file_dump fifo_csv_dumper_958;
    csv_file_dump cstatus_csv_dumper_958;
    df_fifo_monitor fifo_monitor_958;
    df_fifo_intf fifo_intf_959(clock,reset);
    assign fifo_intf_959.rd_en = AESL_inst_myproject.layer2_out_958_U.if_read & AESL_inst_myproject.layer2_out_958_U.if_empty_n;
    assign fifo_intf_959.wr_en = AESL_inst_myproject.layer2_out_958_U.if_write & AESL_inst_myproject.layer2_out_958_U.if_full_n;
    assign fifo_intf_959.fifo_rd_block = 0;
    assign fifo_intf_959.fifo_wr_block = 0;
    assign fifo_intf_959.finish = finish;
    csv_file_dump fifo_csv_dumper_959;
    csv_file_dump cstatus_csv_dumper_959;
    df_fifo_monitor fifo_monitor_959;
    df_fifo_intf fifo_intf_960(clock,reset);
    assign fifo_intf_960.rd_en = AESL_inst_myproject.layer2_out_959_U.if_read & AESL_inst_myproject.layer2_out_959_U.if_empty_n;
    assign fifo_intf_960.wr_en = AESL_inst_myproject.layer2_out_959_U.if_write & AESL_inst_myproject.layer2_out_959_U.if_full_n;
    assign fifo_intf_960.fifo_rd_block = 0;
    assign fifo_intf_960.fifo_wr_block = 0;
    assign fifo_intf_960.finish = finish;
    csv_file_dump fifo_csv_dumper_960;
    csv_file_dump cstatus_csv_dumper_960;
    df_fifo_monitor fifo_monitor_960;
    df_fifo_intf fifo_intf_961(clock,reset);
    assign fifo_intf_961.rd_en = AESL_inst_myproject.layer2_out_960_U.if_read & AESL_inst_myproject.layer2_out_960_U.if_empty_n;
    assign fifo_intf_961.wr_en = AESL_inst_myproject.layer2_out_960_U.if_write & AESL_inst_myproject.layer2_out_960_U.if_full_n;
    assign fifo_intf_961.fifo_rd_block = 0;
    assign fifo_intf_961.fifo_wr_block = 0;
    assign fifo_intf_961.finish = finish;
    csv_file_dump fifo_csv_dumper_961;
    csv_file_dump cstatus_csv_dumper_961;
    df_fifo_monitor fifo_monitor_961;
    df_fifo_intf fifo_intf_962(clock,reset);
    assign fifo_intf_962.rd_en = AESL_inst_myproject.layer2_out_961_U.if_read & AESL_inst_myproject.layer2_out_961_U.if_empty_n;
    assign fifo_intf_962.wr_en = AESL_inst_myproject.layer2_out_961_U.if_write & AESL_inst_myproject.layer2_out_961_U.if_full_n;
    assign fifo_intf_962.fifo_rd_block = 0;
    assign fifo_intf_962.fifo_wr_block = 0;
    assign fifo_intf_962.finish = finish;
    csv_file_dump fifo_csv_dumper_962;
    csv_file_dump cstatus_csv_dumper_962;
    df_fifo_monitor fifo_monitor_962;
    df_fifo_intf fifo_intf_963(clock,reset);
    assign fifo_intf_963.rd_en = AESL_inst_myproject.layer2_out_962_U.if_read & AESL_inst_myproject.layer2_out_962_U.if_empty_n;
    assign fifo_intf_963.wr_en = AESL_inst_myproject.layer2_out_962_U.if_write & AESL_inst_myproject.layer2_out_962_U.if_full_n;
    assign fifo_intf_963.fifo_rd_block = 0;
    assign fifo_intf_963.fifo_wr_block = 0;
    assign fifo_intf_963.finish = finish;
    csv_file_dump fifo_csv_dumper_963;
    csv_file_dump cstatus_csv_dumper_963;
    df_fifo_monitor fifo_monitor_963;
    df_fifo_intf fifo_intf_964(clock,reset);
    assign fifo_intf_964.rd_en = AESL_inst_myproject.layer2_out_963_U.if_read & AESL_inst_myproject.layer2_out_963_U.if_empty_n;
    assign fifo_intf_964.wr_en = AESL_inst_myproject.layer2_out_963_U.if_write & AESL_inst_myproject.layer2_out_963_U.if_full_n;
    assign fifo_intf_964.fifo_rd_block = 0;
    assign fifo_intf_964.fifo_wr_block = 0;
    assign fifo_intf_964.finish = finish;
    csv_file_dump fifo_csv_dumper_964;
    csv_file_dump cstatus_csv_dumper_964;
    df_fifo_monitor fifo_monitor_964;
    df_fifo_intf fifo_intf_965(clock,reset);
    assign fifo_intf_965.rd_en = AESL_inst_myproject.layer2_out_964_U.if_read & AESL_inst_myproject.layer2_out_964_U.if_empty_n;
    assign fifo_intf_965.wr_en = AESL_inst_myproject.layer2_out_964_U.if_write & AESL_inst_myproject.layer2_out_964_U.if_full_n;
    assign fifo_intf_965.fifo_rd_block = 0;
    assign fifo_intf_965.fifo_wr_block = 0;
    assign fifo_intf_965.finish = finish;
    csv_file_dump fifo_csv_dumper_965;
    csv_file_dump cstatus_csv_dumper_965;
    df_fifo_monitor fifo_monitor_965;
    df_fifo_intf fifo_intf_966(clock,reset);
    assign fifo_intf_966.rd_en = AESL_inst_myproject.layer2_out_965_U.if_read & AESL_inst_myproject.layer2_out_965_U.if_empty_n;
    assign fifo_intf_966.wr_en = AESL_inst_myproject.layer2_out_965_U.if_write & AESL_inst_myproject.layer2_out_965_U.if_full_n;
    assign fifo_intf_966.fifo_rd_block = 0;
    assign fifo_intf_966.fifo_wr_block = 0;
    assign fifo_intf_966.finish = finish;
    csv_file_dump fifo_csv_dumper_966;
    csv_file_dump cstatus_csv_dumper_966;
    df_fifo_monitor fifo_monitor_966;
    df_fifo_intf fifo_intf_967(clock,reset);
    assign fifo_intf_967.rd_en = AESL_inst_myproject.layer2_out_966_U.if_read & AESL_inst_myproject.layer2_out_966_U.if_empty_n;
    assign fifo_intf_967.wr_en = AESL_inst_myproject.layer2_out_966_U.if_write & AESL_inst_myproject.layer2_out_966_U.if_full_n;
    assign fifo_intf_967.fifo_rd_block = 0;
    assign fifo_intf_967.fifo_wr_block = 0;
    assign fifo_intf_967.finish = finish;
    csv_file_dump fifo_csv_dumper_967;
    csv_file_dump cstatus_csv_dumper_967;
    df_fifo_monitor fifo_monitor_967;
    df_fifo_intf fifo_intf_968(clock,reset);
    assign fifo_intf_968.rd_en = AESL_inst_myproject.layer2_out_967_U.if_read & AESL_inst_myproject.layer2_out_967_U.if_empty_n;
    assign fifo_intf_968.wr_en = AESL_inst_myproject.layer2_out_967_U.if_write & AESL_inst_myproject.layer2_out_967_U.if_full_n;
    assign fifo_intf_968.fifo_rd_block = 0;
    assign fifo_intf_968.fifo_wr_block = 0;
    assign fifo_intf_968.finish = finish;
    csv_file_dump fifo_csv_dumper_968;
    csv_file_dump cstatus_csv_dumper_968;
    df_fifo_monitor fifo_monitor_968;
    df_fifo_intf fifo_intf_969(clock,reset);
    assign fifo_intf_969.rd_en = AESL_inst_myproject.layer2_out_968_U.if_read & AESL_inst_myproject.layer2_out_968_U.if_empty_n;
    assign fifo_intf_969.wr_en = AESL_inst_myproject.layer2_out_968_U.if_write & AESL_inst_myproject.layer2_out_968_U.if_full_n;
    assign fifo_intf_969.fifo_rd_block = 0;
    assign fifo_intf_969.fifo_wr_block = 0;
    assign fifo_intf_969.finish = finish;
    csv_file_dump fifo_csv_dumper_969;
    csv_file_dump cstatus_csv_dumper_969;
    df_fifo_monitor fifo_monitor_969;
    df_fifo_intf fifo_intf_970(clock,reset);
    assign fifo_intf_970.rd_en = AESL_inst_myproject.layer2_out_969_U.if_read & AESL_inst_myproject.layer2_out_969_U.if_empty_n;
    assign fifo_intf_970.wr_en = AESL_inst_myproject.layer2_out_969_U.if_write & AESL_inst_myproject.layer2_out_969_U.if_full_n;
    assign fifo_intf_970.fifo_rd_block = 0;
    assign fifo_intf_970.fifo_wr_block = 0;
    assign fifo_intf_970.finish = finish;
    csv_file_dump fifo_csv_dumper_970;
    csv_file_dump cstatus_csv_dumper_970;
    df_fifo_monitor fifo_monitor_970;
    df_fifo_intf fifo_intf_971(clock,reset);
    assign fifo_intf_971.rd_en = AESL_inst_myproject.layer2_out_970_U.if_read & AESL_inst_myproject.layer2_out_970_U.if_empty_n;
    assign fifo_intf_971.wr_en = AESL_inst_myproject.layer2_out_970_U.if_write & AESL_inst_myproject.layer2_out_970_U.if_full_n;
    assign fifo_intf_971.fifo_rd_block = 0;
    assign fifo_intf_971.fifo_wr_block = 0;
    assign fifo_intf_971.finish = finish;
    csv_file_dump fifo_csv_dumper_971;
    csv_file_dump cstatus_csv_dumper_971;
    df_fifo_monitor fifo_monitor_971;
    df_fifo_intf fifo_intf_972(clock,reset);
    assign fifo_intf_972.rd_en = AESL_inst_myproject.layer2_out_971_U.if_read & AESL_inst_myproject.layer2_out_971_U.if_empty_n;
    assign fifo_intf_972.wr_en = AESL_inst_myproject.layer2_out_971_U.if_write & AESL_inst_myproject.layer2_out_971_U.if_full_n;
    assign fifo_intf_972.fifo_rd_block = 0;
    assign fifo_intf_972.fifo_wr_block = 0;
    assign fifo_intf_972.finish = finish;
    csv_file_dump fifo_csv_dumper_972;
    csv_file_dump cstatus_csv_dumper_972;
    df_fifo_monitor fifo_monitor_972;
    df_fifo_intf fifo_intf_973(clock,reset);
    assign fifo_intf_973.rd_en = AESL_inst_myproject.layer2_out_972_U.if_read & AESL_inst_myproject.layer2_out_972_U.if_empty_n;
    assign fifo_intf_973.wr_en = AESL_inst_myproject.layer2_out_972_U.if_write & AESL_inst_myproject.layer2_out_972_U.if_full_n;
    assign fifo_intf_973.fifo_rd_block = 0;
    assign fifo_intf_973.fifo_wr_block = 0;
    assign fifo_intf_973.finish = finish;
    csv_file_dump fifo_csv_dumper_973;
    csv_file_dump cstatus_csv_dumper_973;
    df_fifo_monitor fifo_monitor_973;
    df_fifo_intf fifo_intf_974(clock,reset);
    assign fifo_intf_974.rd_en = AESL_inst_myproject.layer2_out_973_U.if_read & AESL_inst_myproject.layer2_out_973_U.if_empty_n;
    assign fifo_intf_974.wr_en = AESL_inst_myproject.layer2_out_973_U.if_write & AESL_inst_myproject.layer2_out_973_U.if_full_n;
    assign fifo_intf_974.fifo_rd_block = 0;
    assign fifo_intf_974.fifo_wr_block = 0;
    assign fifo_intf_974.finish = finish;
    csv_file_dump fifo_csv_dumper_974;
    csv_file_dump cstatus_csv_dumper_974;
    df_fifo_monitor fifo_monitor_974;
    df_fifo_intf fifo_intf_975(clock,reset);
    assign fifo_intf_975.rd_en = AESL_inst_myproject.layer2_out_974_U.if_read & AESL_inst_myproject.layer2_out_974_U.if_empty_n;
    assign fifo_intf_975.wr_en = AESL_inst_myproject.layer2_out_974_U.if_write & AESL_inst_myproject.layer2_out_974_U.if_full_n;
    assign fifo_intf_975.fifo_rd_block = 0;
    assign fifo_intf_975.fifo_wr_block = 0;
    assign fifo_intf_975.finish = finish;
    csv_file_dump fifo_csv_dumper_975;
    csv_file_dump cstatus_csv_dumper_975;
    df_fifo_monitor fifo_monitor_975;
    df_fifo_intf fifo_intf_976(clock,reset);
    assign fifo_intf_976.rd_en = AESL_inst_myproject.layer2_out_975_U.if_read & AESL_inst_myproject.layer2_out_975_U.if_empty_n;
    assign fifo_intf_976.wr_en = AESL_inst_myproject.layer2_out_975_U.if_write & AESL_inst_myproject.layer2_out_975_U.if_full_n;
    assign fifo_intf_976.fifo_rd_block = 0;
    assign fifo_intf_976.fifo_wr_block = 0;
    assign fifo_intf_976.finish = finish;
    csv_file_dump fifo_csv_dumper_976;
    csv_file_dump cstatus_csv_dumper_976;
    df_fifo_monitor fifo_monitor_976;
    df_fifo_intf fifo_intf_977(clock,reset);
    assign fifo_intf_977.rd_en = AESL_inst_myproject.layer2_out_976_U.if_read & AESL_inst_myproject.layer2_out_976_U.if_empty_n;
    assign fifo_intf_977.wr_en = AESL_inst_myproject.layer2_out_976_U.if_write & AESL_inst_myproject.layer2_out_976_U.if_full_n;
    assign fifo_intf_977.fifo_rd_block = 0;
    assign fifo_intf_977.fifo_wr_block = 0;
    assign fifo_intf_977.finish = finish;
    csv_file_dump fifo_csv_dumper_977;
    csv_file_dump cstatus_csv_dumper_977;
    df_fifo_monitor fifo_monitor_977;
    df_fifo_intf fifo_intf_978(clock,reset);
    assign fifo_intf_978.rd_en = AESL_inst_myproject.layer2_out_977_U.if_read & AESL_inst_myproject.layer2_out_977_U.if_empty_n;
    assign fifo_intf_978.wr_en = AESL_inst_myproject.layer2_out_977_U.if_write & AESL_inst_myproject.layer2_out_977_U.if_full_n;
    assign fifo_intf_978.fifo_rd_block = 0;
    assign fifo_intf_978.fifo_wr_block = 0;
    assign fifo_intf_978.finish = finish;
    csv_file_dump fifo_csv_dumper_978;
    csv_file_dump cstatus_csv_dumper_978;
    df_fifo_monitor fifo_monitor_978;
    df_fifo_intf fifo_intf_979(clock,reset);
    assign fifo_intf_979.rd_en = AESL_inst_myproject.layer2_out_978_U.if_read & AESL_inst_myproject.layer2_out_978_U.if_empty_n;
    assign fifo_intf_979.wr_en = AESL_inst_myproject.layer2_out_978_U.if_write & AESL_inst_myproject.layer2_out_978_U.if_full_n;
    assign fifo_intf_979.fifo_rd_block = 0;
    assign fifo_intf_979.fifo_wr_block = 0;
    assign fifo_intf_979.finish = finish;
    csv_file_dump fifo_csv_dumper_979;
    csv_file_dump cstatus_csv_dumper_979;
    df_fifo_monitor fifo_monitor_979;
    df_fifo_intf fifo_intf_980(clock,reset);
    assign fifo_intf_980.rd_en = AESL_inst_myproject.layer2_out_979_U.if_read & AESL_inst_myproject.layer2_out_979_U.if_empty_n;
    assign fifo_intf_980.wr_en = AESL_inst_myproject.layer2_out_979_U.if_write & AESL_inst_myproject.layer2_out_979_U.if_full_n;
    assign fifo_intf_980.fifo_rd_block = 0;
    assign fifo_intf_980.fifo_wr_block = 0;
    assign fifo_intf_980.finish = finish;
    csv_file_dump fifo_csv_dumper_980;
    csv_file_dump cstatus_csv_dumper_980;
    df_fifo_monitor fifo_monitor_980;
    df_fifo_intf fifo_intf_981(clock,reset);
    assign fifo_intf_981.rd_en = AESL_inst_myproject.layer2_out_980_U.if_read & AESL_inst_myproject.layer2_out_980_U.if_empty_n;
    assign fifo_intf_981.wr_en = AESL_inst_myproject.layer2_out_980_U.if_write & AESL_inst_myproject.layer2_out_980_U.if_full_n;
    assign fifo_intf_981.fifo_rd_block = 0;
    assign fifo_intf_981.fifo_wr_block = 0;
    assign fifo_intf_981.finish = finish;
    csv_file_dump fifo_csv_dumper_981;
    csv_file_dump cstatus_csv_dumper_981;
    df_fifo_monitor fifo_monitor_981;
    df_fifo_intf fifo_intf_982(clock,reset);
    assign fifo_intf_982.rd_en = AESL_inst_myproject.layer2_out_981_U.if_read & AESL_inst_myproject.layer2_out_981_U.if_empty_n;
    assign fifo_intf_982.wr_en = AESL_inst_myproject.layer2_out_981_U.if_write & AESL_inst_myproject.layer2_out_981_U.if_full_n;
    assign fifo_intf_982.fifo_rd_block = 0;
    assign fifo_intf_982.fifo_wr_block = 0;
    assign fifo_intf_982.finish = finish;
    csv_file_dump fifo_csv_dumper_982;
    csv_file_dump cstatus_csv_dumper_982;
    df_fifo_monitor fifo_monitor_982;
    df_fifo_intf fifo_intf_983(clock,reset);
    assign fifo_intf_983.rd_en = AESL_inst_myproject.layer2_out_982_U.if_read & AESL_inst_myproject.layer2_out_982_U.if_empty_n;
    assign fifo_intf_983.wr_en = AESL_inst_myproject.layer2_out_982_U.if_write & AESL_inst_myproject.layer2_out_982_U.if_full_n;
    assign fifo_intf_983.fifo_rd_block = 0;
    assign fifo_intf_983.fifo_wr_block = 0;
    assign fifo_intf_983.finish = finish;
    csv_file_dump fifo_csv_dumper_983;
    csv_file_dump cstatus_csv_dumper_983;
    df_fifo_monitor fifo_monitor_983;
    df_fifo_intf fifo_intf_984(clock,reset);
    assign fifo_intf_984.rd_en = AESL_inst_myproject.layer2_out_983_U.if_read & AESL_inst_myproject.layer2_out_983_U.if_empty_n;
    assign fifo_intf_984.wr_en = AESL_inst_myproject.layer2_out_983_U.if_write & AESL_inst_myproject.layer2_out_983_U.if_full_n;
    assign fifo_intf_984.fifo_rd_block = 0;
    assign fifo_intf_984.fifo_wr_block = 0;
    assign fifo_intf_984.finish = finish;
    csv_file_dump fifo_csv_dumper_984;
    csv_file_dump cstatus_csv_dumper_984;
    df_fifo_monitor fifo_monitor_984;
    df_fifo_intf fifo_intf_985(clock,reset);
    assign fifo_intf_985.rd_en = AESL_inst_myproject.layer2_out_984_U.if_read & AESL_inst_myproject.layer2_out_984_U.if_empty_n;
    assign fifo_intf_985.wr_en = AESL_inst_myproject.layer2_out_984_U.if_write & AESL_inst_myproject.layer2_out_984_U.if_full_n;
    assign fifo_intf_985.fifo_rd_block = 0;
    assign fifo_intf_985.fifo_wr_block = 0;
    assign fifo_intf_985.finish = finish;
    csv_file_dump fifo_csv_dumper_985;
    csv_file_dump cstatus_csv_dumper_985;
    df_fifo_monitor fifo_monitor_985;
    df_fifo_intf fifo_intf_986(clock,reset);
    assign fifo_intf_986.rd_en = AESL_inst_myproject.layer2_out_985_U.if_read & AESL_inst_myproject.layer2_out_985_U.if_empty_n;
    assign fifo_intf_986.wr_en = AESL_inst_myproject.layer2_out_985_U.if_write & AESL_inst_myproject.layer2_out_985_U.if_full_n;
    assign fifo_intf_986.fifo_rd_block = 0;
    assign fifo_intf_986.fifo_wr_block = 0;
    assign fifo_intf_986.finish = finish;
    csv_file_dump fifo_csv_dumper_986;
    csv_file_dump cstatus_csv_dumper_986;
    df_fifo_monitor fifo_monitor_986;
    df_fifo_intf fifo_intf_987(clock,reset);
    assign fifo_intf_987.rd_en = AESL_inst_myproject.layer2_out_986_U.if_read & AESL_inst_myproject.layer2_out_986_U.if_empty_n;
    assign fifo_intf_987.wr_en = AESL_inst_myproject.layer2_out_986_U.if_write & AESL_inst_myproject.layer2_out_986_U.if_full_n;
    assign fifo_intf_987.fifo_rd_block = 0;
    assign fifo_intf_987.fifo_wr_block = 0;
    assign fifo_intf_987.finish = finish;
    csv_file_dump fifo_csv_dumper_987;
    csv_file_dump cstatus_csv_dumper_987;
    df_fifo_monitor fifo_monitor_987;
    df_fifo_intf fifo_intf_988(clock,reset);
    assign fifo_intf_988.rd_en = AESL_inst_myproject.layer2_out_987_U.if_read & AESL_inst_myproject.layer2_out_987_U.if_empty_n;
    assign fifo_intf_988.wr_en = AESL_inst_myproject.layer2_out_987_U.if_write & AESL_inst_myproject.layer2_out_987_U.if_full_n;
    assign fifo_intf_988.fifo_rd_block = 0;
    assign fifo_intf_988.fifo_wr_block = 0;
    assign fifo_intf_988.finish = finish;
    csv_file_dump fifo_csv_dumper_988;
    csv_file_dump cstatus_csv_dumper_988;
    df_fifo_monitor fifo_monitor_988;
    df_fifo_intf fifo_intf_989(clock,reset);
    assign fifo_intf_989.rd_en = AESL_inst_myproject.layer2_out_988_U.if_read & AESL_inst_myproject.layer2_out_988_U.if_empty_n;
    assign fifo_intf_989.wr_en = AESL_inst_myproject.layer2_out_988_U.if_write & AESL_inst_myproject.layer2_out_988_U.if_full_n;
    assign fifo_intf_989.fifo_rd_block = 0;
    assign fifo_intf_989.fifo_wr_block = 0;
    assign fifo_intf_989.finish = finish;
    csv_file_dump fifo_csv_dumper_989;
    csv_file_dump cstatus_csv_dumper_989;
    df_fifo_monitor fifo_monitor_989;
    df_fifo_intf fifo_intf_990(clock,reset);
    assign fifo_intf_990.rd_en = AESL_inst_myproject.layer2_out_989_U.if_read & AESL_inst_myproject.layer2_out_989_U.if_empty_n;
    assign fifo_intf_990.wr_en = AESL_inst_myproject.layer2_out_989_U.if_write & AESL_inst_myproject.layer2_out_989_U.if_full_n;
    assign fifo_intf_990.fifo_rd_block = 0;
    assign fifo_intf_990.fifo_wr_block = 0;
    assign fifo_intf_990.finish = finish;
    csv_file_dump fifo_csv_dumper_990;
    csv_file_dump cstatus_csv_dumper_990;
    df_fifo_monitor fifo_monitor_990;
    df_fifo_intf fifo_intf_991(clock,reset);
    assign fifo_intf_991.rd_en = AESL_inst_myproject.layer2_out_990_U.if_read & AESL_inst_myproject.layer2_out_990_U.if_empty_n;
    assign fifo_intf_991.wr_en = AESL_inst_myproject.layer2_out_990_U.if_write & AESL_inst_myproject.layer2_out_990_U.if_full_n;
    assign fifo_intf_991.fifo_rd_block = 0;
    assign fifo_intf_991.fifo_wr_block = 0;
    assign fifo_intf_991.finish = finish;
    csv_file_dump fifo_csv_dumper_991;
    csv_file_dump cstatus_csv_dumper_991;
    df_fifo_monitor fifo_monitor_991;
    df_fifo_intf fifo_intf_992(clock,reset);
    assign fifo_intf_992.rd_en = AESL_inst_myproject.layer2_out_991_U.if_read & AESL_inst_myproject.layer2_out_991_U.if_empty_n;
    assign fifo_intf_992.wr_en = AESL_inst_myproject.layer2_out_991_U.if_write & AESL_inst_myproject.layer2_out_991_U.if_full_n;
    assign fifo_intf_992.fifo_rd_block = 0;
    assign fifo_intf_992.fifo_wr_block = 0;
    assign fifo_intf_992.finish = finish;
    csv_file_dump fifo_csv_dumper_992;
    csv_file_dump cstatus_csv_dumper_992;
    df_fifo_monitor fifo_monitor_992;
    df_fifo_intf fifo_intf_993(clock,reset);
    assign fifo_intf_993.rd_en = AESL_inst_myproject.layer2_out_992_U.if_read & AESL_inst_myproject.layer2_out_992_U.if_empty_n;
    assign fifo_intf_993.wr_en = AESL_inst_myproject.layer2_out_992_U.if_write & AESL_inst_myproject.layer2_out_992_U.if_full_n;
    assign fifo_intf_993.fifo_rd_block = 0;
    assign fifo_intf_993.fifo_wr_block = 0;
    assign fifo_intf_993.finish = finish;
    csv_file_dump fifo_csv_dumper_993;
    csv_file_dump cstatus_csv_dumper_993;
    df_fifo_monitor fifo_monitor_993;
    df_fifo_intf fifo_intf_994(clock,reset);
    assign fifo_intf_994.rd_en = AESL_inst_myproject.layer2_out_993_U.if_read & AESL_inst_myproject.layer2_out_993_U.if_empty_n;
    assign fifo_intf_994.wr_en = AESL_inst_myproject.layer2_out_993_U.if_write & AESL_inst_myproject.layer2_out_993_U.if_full_n;
    assign fifo_intf_994.fifo_rd_block = 0;
    assign fifo_intf_994.fifo_wr_block = 0;
    assign fifo_intf_994.finish = finish;
    csv_file_dump fifo_csv_dumper_994;
    csv_file_dump cstatus_csv_dumper_994;
    df_fifo_monitor fifo_monitor_994;
    df_fifo_intf fifo_intf_995(clock,reset);
    assign fifo_intf_995.rd_en = AESL_inst_myproject.layer2_out_994_U.if_read & AESL_inst_myproject.layer2_out_994_U.if_empty_n;
    assign fifo_intf_995.wr_en = AESL_inst_myproject.layer2_out_994_U.if_write & AESL_inst_myproject.layer2_out_994_U.if_full_n;
    assign fifo_intf_995.fifo_rd_block = 0;
    assign fifo_intf_995.fifo_wr_block = 0;
    assign fifo_intf_995.finish = finish;
    csv_file_dump fifo_csv_dumper_995;
    csv_file_dump cstatus_csv_dumper_995;
    df_fifo_monitor fifo_monitor_995;
    df_fifo_intf fifo_intf_996(clock,reset);
    assign fifo_intf_996.rd_en = AESL_inst_myproject.layer2_out_995_U.if_read & AESL_inst_myproject.layer2_out_995_U.if_empty_n;
    assign fifo_intf_996.wr_en = AESL_inst_myproject.layer2_out_995_U.if_write & AESL_inst_myproject.layer2_out_995_U.if_full_n;
    assign fifo_intf_996.fifo_rd_block = 0;
    assign fifo_intf_996.fifo_wr_block = 0;
    assign fifo_intf_996.finish = finish;
    csv_file_dump fifo_csv_dumper_996;
    csv_file_dump cstatus_csv_dumper_996;
    df_fifo_monitor fifo_monitor_996;
    df_fifo_intf fifo_intf_997(clock,reset);
    assign fifo_intf_997.rd_en = AESL_inst_myproject.layer2_out_996_U.if_read & AESL_inst_myproject.layer2_out_996_U.if_empty_n;
    assign fifo_intf_997.wr_en = AESL_inst_myproject.layer2_out_996_U.if_write & AESL_inst_myproject.layer2_out_996_U.if_full_n;
    assign fifo_intf_997.fifo_rd_block = 0;
    assign fifo_intf_997.fifo_wr_block = 0;
    assign fifo_intf_997.finish = finish;
    csv_file_dump fifo_csv_dumper_997;
    csv_file_dump cstatus_csv_dumper_997;
    df_fifo_monitor fifo_monitor_997;
    df_fifo_intf fifo_intf_998(clock,reset);
    assign fifo_intf_998.rd_en = AESL_inst_myproject.layer2_out_997_U.if_read & AESL_inst_myproject.layer2_out_997_U.if_empty_n;
    assign fifo_intf_998.wr_en = AESL_inst_myproject.layer2_out_997_U.if_write & AESL_inst_myproject.layer2_out_997_U.if_full_n;
    assign fifo_intf_998.fifo_rd_block = 0;
    assign fifo_intf_998.fifo_wr_block = 0;
    assign fifo_intf_998.finish = finish;
    csv_file_dump fifo_csv_dumper_998;
    csv_file_dump cstatus_csv_dumper_998;
    df_fifo_monitor fifo_monitor_998;
    df_fifo_intf fifo_intf_999(clock,reset);
    assign fifo_intf_999.rd_en = AESL_inst_myproject.layer2_out_998_U.if_read & AESL_inst_myproject.layer2_out_998_U.if_empty_n;
    assign fifo_intf_999.wr_en = AESL_inst_myproject.layer2_out_998_U.if_write & AESL_inst_myproject.layer2_out_998_U.if_full_n;
    assign fifo_intf_999.fifo_rd_block = 0;
    assign fifo_intf_999.fifo_wr_block = 0;
    assign fifo_intf_999.finish = finish;
    csv_file_dump fifo_csv_dumper_999;
    csv_file_dump cstatus_csv_dumper_999;
    df_fifo_monitor fifo_monitor_999;
    df_fifo_intf fifo_intf_1000(clock,reset);
    assign fifo_intf_1000.rd_en = AESL_inst_myproject.layer2_out_999_U.if_read & AESL_inst_myproject.layer2_out_999_U.if_empty_n;
    assign fifo_intf_1000.wr_en = AESL_inst_myproject.layer2_out_999_U.if_write & AESL_inst_myproject.layer2_out_999_U.if_full_n;
    assign fifo_intf_1000.fifo_rd_block = 0;
    assign fifo_intf_1000.fifo_wr_block = 0;
    assign fifo_intf_1000.finish = finish;
    csv_file_dump fifo_csv_dumper_1000;
    csv_file_dump cstatus_csv_dumper_1000;
    df_fifo_monitor fifo_monitor_1000;
    df_fifo_intf fifo_intf_1001(clock,reset);
    assign fifo_intf_1001.rd_en = AESL_inst_myproject.layer2_out_1000_U.if_read & AESL_inst_myproject.layer2_out_1000_U.if_empty_n;
    assign fifo_intf_1001.wr_en = AESL_inst_myproject.layer2_out_1000_U.if_write & AESL_inst_myproject.layer2_out_1000_U.if_full_n;
    assign fifo_intf_1001.fifo_rd_block = 0;
    assign fifo_intf_1001.fifo_wr_block = 0;
    assign fifo_intf_1001.finish = finish;
    csv_file_dump fifo_csv_dumper_1001;
    csv_file_dump cstatus_csv_dumper_1001;
    df_fifo_monitor fifo_monitor_1001;
    df_fifo_intf fifo_intf_1002(clock,reset);
    assign fifo_intf_1002.rd_en = AESL_inst_myproject.layer2_out_1001_U.if_read & AESL_inst_myproject.layer2_out_1001_U.if_empty_n;
    assign fifo_intf_1002.wr_en = AESL_inst_myproject.layer2_out_1001_U.if_write & AESL_inst_myproject.layer2_out_1001_U.if_full_n;
    assign fifo_intf_1002.fifo_rd_block = 0;
    assign fifo_intf_1002.fifo_wr_block = 0;
    assign fifo_intf_1002.finish = finish;
    csv_file_dump fifo_csv_dumper_1002;
    csv_file_dump cstatus_csv_dumper_1002;
    df_fifo_monitor fifo_monitor_1002;
    df_fifo_intf fifo_intf_1003(clock,reset);
    assign fifo_intf_1003.rd_en = AESL_inst_myproject.layer2_out_1002_U.if_read & AESL_inst_myproject.layer2_out_1002_U.if_empty_n;
    assign fifo_intf_1003.wr_en = AESL_inst_myproject.layer2_out_1002_U.if_write & AESL_inst_myproject.layer2_out_1002_U.if_full_n;
    assign fifo_intf_1003.fifo_rd_block = 0;
    assign fifo_intf_1003.fifo_wr_block = 0;
    assign fifo_intf_1003.finish = finish;
    csv_file_dump fifo_csv_dumper_1003;
    csv_file_dump cstatus_csv_dumper_1003;
    df_fifo_monitor fifo_monitor_1003;
    df_fifo_intf fifo_intf_1004(clock,reset);
    assign fifo_intf_1004.rd_en = AESL_inst_myproject.layer2_out_1003_U.if_read & AESL_inst_myproject.layer2_out_1003_U.if_empty_n;
    assign fifo_intf_1004.wr_en = AESL_inst_myproject.layer2_out_1003_U.if_write & AESL_inst_myproject.layer2_out_1003_U.if_full_n;
    assign fifo_intf_1004.fifo_rd_block = 0;
    assign fifo_intf_1004.fifo_wr_block = 0;
    assign fifo_intf_1004.finish = finish;
    csv_file_dump fifo_csv_dumper_1004;
    csv_file_dump cstatus_csv_dumper_1004;
    df_fifo_monitor fifo_monitor_1004;
    df_fifo_intf fifo_intf_1005(clock,reset);
    assign fifo_intf_1005.rd_en = AESL_inst_myproject.layer2_out_1004_U.if_read & AESL_inst_myproject.layer2_out_1004_U.if_empty_n;
    assign fifo_intf_1005.wr_en = AESL_inst_myproject.layer2_out_1004_U.if_write & AESL_inst_myproject.layer2_out_1004_U.if_full_n;
    assign fifo_intf_1005.fifo_rd_block = 0;
    assign fifo_intf_1005.fifo_wr_block = 0;
    assign fifo_intf_1005.finish = finish;
    csv_file_dump fifo_csv_dumper_1005;
    csv_file_dump cstatus_csv_dumper_1005;
    df_fifo_monitor fifo_monitor_1005;
    df_fifo_intf fifo_intf_1006(clock,reset);
    assign fifo_intf_1006.rd_en = AESL_inst_myproject.layer2_out_1005_U.if_read & AESL_inst_myproject.layer2_out_1005_U.if_empty_n;
    assign fifo_intf_1006.wr_en = AESL_inst_myproject.layer2_out_1005_U.if_write & AESL_inst_myproject.layer2_out_1005_U.if_full_n;
    assign fifo_intf_1006.fifo_rd_block = 0;
    assign fifo_intf_1006.fifo_wr_block = 0;
    assign fifo_intf_1006.finish = finish;
    csv_file_dump fifo_csv_dumper_1006;
    csv_file_dump cstatus_csv_dumper_1006;
    df_fifo_monitor fifo_monitor_1006;
    df_fifo_intf fifo_intf_1007(clock,reset);
    assign fifo_intf_1007.rd_en = AESL_inst_myproject.layer2_out_1006_U.if_read & AESL_inst_myproject.layer2_out_1006_U.if_empty_n;
    assign fifo_intf_1007.wr_en = AESL_inst_myproject.layer2_out_1006_U.if_write & AESL_inst_myproject.layer2_out_1006_U.if_full_n;
    assign fifo_intf_1007.fifo_rd_block = 0;
    assign fifo_intf_1007.fifo_wr_block = 0;
    assign fifo_intf_1007.finish = finish;
    csv_file_dump fifo_csv_dumper_1007;
    csv_file_dump cstatus_csv_dumper_1007;
    df_fifo_monitor fifo_monitor_1007;
    df_fifo_intf fifo_intf_1008(clock,reset);
    assign fifo_intf_1008.rd_en = AESL_inst_myproject.layer2_out_1007_U.if_read & AESL_inst_myproject.layer2_out_1007_U.if_empty_n;
    assign fifo_intf_1008.wr_en = AESL_inst_myproject.layer2_out_1007_U.if_write & AESL_inst_myproject.layer2_out_1007_U.if_full_n;
    assign fifo_intf_1008.fifo_rd_block = 0;
    assign fifo_intf_1008.fifo_wr_block = 0;
    assign fifo_intf_1008.finish = finish;
    csv_file_dump fifo_csv_dumper_1008;
    csv_file_dump cstatus_csv_dumper_1008;
    df_fifo_monitor fifo_monitor_1008;
    df_fifo_intf fifo_intf_1009(clock,reset);
    assign fifo_intf_1009.rd_en = AESL_inst_myproject.layer2_out_1008_U.if_read & AESL_inst_myproject.layer2_out_1008_U.if_empty_n;
    assign fifo_intf_1009.wr_en = AESL_inst_myproject.layer2_out_1008_U.if_write & AESL_inst_myproject.layer2_out_1008_U.if_full_n;
    assign fifo_intf_1009.fifo_rd_block = 0;
    assign fifo_intf_1009.fifo_wr_block = 0;
    assign fifo_intf_1009.finish = finish;
    csv_file_dump fifo_csv_dumper_1009;
    csv_file_dump cstatus_csv_dumper_1009;
    df_fifo_monitor fifo_monitor_1009;
    df_fifo_intf fifo_intf_1010(clock,reset);
    assign fifo_intf_1010.rd_en = AESL_inst_myproject.layer2_out_1009_U.if_read & AESL_inst_myproject.layer2_out_1009_U.if_empty_n;
    assign fifo_intf_1010.wr_en = AESL_inst_myproject.layer2_out_1009_U.if_write & AESL_inst_myproject.layer2_out_1009_U.if_full_n;
    assign fifo_intf_1010.fifo_rd_block = 0;
    assign fifo_intf_1010.fifo_wr_block = 0;
    assign fifo_intf_1010.finish = finish;
    csv_file_dump fifo_csv_dumper_1010;
    csv_file_dump cstatus_csv_dumper_1010;
    df_fifo_monitor fifo_monitor_1010;
    df_fifo_intf fifo_intf_1011(clock,reset);
    assign fifo_intf_1011.rd_en = AESL_inst_myproject.layer2_out_1010_U.if_read & AESL_inst_myproject.layer2_out_1010_U.if_empty_n;
    assign fifo_intf_1011.wr_en = AESL_inst_myproject.layer2_out_1010_U.if_write & AESL_inst_myproject.layer2_out_1010_U.if_full_n;
    assign fifo_intf_1011.fifo_rd_block = 0;
    assign fifo_intf_1011.fifo_wr_block = 0;
    assign fifo_intf_1011.finish = finish;
    csv_file_dump fifo_csv_dumper_1011;
    csv_file_dump cstatus_csv_dumper_1011;
    df_fifo_monitor fifo_monitor_1011;
    df_fifo_intf fifo_intf_1012(clock,reset);
    assign fifo_intf_1012.rd_en = AESL_inst_myproject.layer2_out_1011_U.if_read & AESL_inst_myproject.layer2_out_1011_U.if_empty_n;
    assign fifo_intf_1012.wr_en = AESL_inst_myproject.layer2_out_1011_U.if_write & AESL_inst_myproject.layer2_out_1011_U.if_full_n;
    assign fifo_intf_1012.fifo_rd_block = 0;
    assign fifo_intf_1012.fifo_wr_block = 0;
    assign fifo_intf_1012.finish = finish;
    csv_file_dump fifo_csv_dumper_1012;
    csv_file_dump cstatus_csv_dumper_1012;
    df_fifo_monitor fifo_monitor_1012;
    df_fifo_intf fifo_intf_1013(clock,reset);
    assign fifo_intf_1013.rd_en = AESL_inst_myproject.layer2_out_1012_U.if_read & AESL_inst_myproject.layer2_out_1012_U.if_empty_n;
    assign fifo_intf_1013.wr_en = AESL_inst_myproject.layer2_out_1012_U.if_write & AESL_inst_myproject.layer2_out_1012_U.if_full_n;
    assign fifo_intf_1013.fifo_rd_block = 0;
    assign fifo_intf_1013.fifo_wr_block = 0;
    assign fifo_intf_1013.finish = finish;
    csv_file_dump fifo_csv_dumper_1013;
    csv_file_dump cstatus_csv_dumper_1013;
    df_fifo_monitor fifo_monitor_1013;
    df_fifo_intf fifo_intf_1014(clock,reset);
    assign fifo_intf_1014.rd_en = AESL_inst_myproject.layer2_out_1013_U.if_read & AESL_inst_myproject.layer2_out_1013_U.if_empty_n;
    assign fifo_intf_1014.wr_en = AESL_inst_myproject.layer2_out_1013_U.if_write & AESL_inst_myproject.layer2_out_1013_U.if_full_n;
    assign fifo_intf_1014.fifo_rd_block = 0;
    assign fifo_intf_1014.fifo_wr_block = 0;
    assign fifo_intf_1014.finish = finish;
    csv_file_dump fifo_csv_dumper_1014;
    csv_file_dump cstatus_csv_dumper_1014;
    df_fifo_monitor fifo_monitor_1014;
    df_fifo_intf fifo_intf_1015(clock,reset);
    assign fifo_intf_1015.rd_en = AESL_inst_myproject.layer2_out_1014_U.if_read & AESL_inst_myproject.layer2_out_1014_U.if_empty_n;
    assign fifo_intf_1015.wr_en = AESL_inst_myproject.layer2_out_1014_U.if_write & AESL_inst_myproject.layer2_out_1014_U.if_full_n;
    assign fifo_intf_1015.fifo_rd_block = 0;
    assign fifo_intf_1015.fifo_wr_block = 0;
    assign fifo_intf_1015.finish = finish;
    csv_file_dump fifo_csv_dumper_1015;
    csv_file_dump cstatus_csv_dumper_1015;
    df_fifo_monitor fifo_monitor_1015;
    df_fifo_intf fifo_intf_1016(clock,reset);
    assign fifo_intf_1016.rd_en = AESL_inst_myproject.layer2_out_1015_U.if_read & AESL_inst_myproject.layer2_out_1015_U.if_empty_n;
    assign fifo_intf_1016.wr_en = AESL_inst_myproject.layer2_out_1015_U.if_write & AESL_inst_myproject.layer2_out_1015_U.if_full_n;
    assign fifo_intf_1016.fifo_rd_block = 0;
    assign fifo_intf_1016.fifo_wr_block = 0;
    assign fifo_intf_1016.finish = finish;
    csv_file_dump fifo_csv_dumper_1016;
    csv_file_dump cstatus_csv_dumper_1016;
    df_fifo_monitor fifo_monitor_1016;
    df_fifo_intf fifo_intf_1017(clock,reset);
    assign fifo_intf_1017.rd_en = AESL_inst_myproject.layer2_out_1016_U.if_read & AESL_inst_myproject.layer2_out_1016_U.if_empty_n;
    assign fifo_intf_1017.wr_en = AESL_inst_myproject.layer2_out_1016_U.if_write & AESL_inst_myproject.layer2_out_1016_U.if_full_n;
    assign fifo_intf_1017.fifo_rd_block = 0;
    assign fifo_intf_1017.fifo_wr_block = 0;
    assign fifo_intf_1017.finish = finish;
    csv_file_dump fifo_csv_dumper_1017;
    csv_file_dump cstatus_csv_dumper_1017;
    df_fifo_monitor fifo_monitor_1017;
    df_fifo_intf fifo_intf_1018(clock,reset);
    assign fifo_intf_1018.rd_en = AESL_inst_myproject.layer2_out_1017_U.if_read & AESL_inst_myproject.layer2_out_1017_U.if_empty_n;
    assign fifo_intf_1018.wr_en = AESL_inst_myproject.layer2_out_1017_U.if_write & AESL_inst_myproject.layer2_out_1017_U.if_full_n;
    assign fifo_intf_1018.fifo_rd_block = 0;
    assign fifo_intf_1018.fifo_wr_block = 0;
    assign fifo_intf_1018.finish = finish;
    csv_file_dump fifo_csv_dumper_1018;
    csv_file_dump cstatus_csv_dumper_1018;
    df_fifo_monitor fifo_monitor_1018;
    df_fifo_intf fifo_intf_1019(clock,reset);
    assign fifo_intf_1019.rd_en = AESL_inst_myproject.layer2_out_1018_U.if_read & AESL_inst_myproject.layer2_out_1018_U.if_empty_n;
    assign fifo_intf_1019.wr_en = AESL_inst_myproject.layer2_out_1018_U.if_write & AESL_inst_myproject.layer2_out_1018_U.if_full_n;
    assign fifo_intf_1019.fifo_rd_block = 0;
    assign fifo_intf_1019.fifo_wr_block = 0;
    assign fifo_intf_1019.finish = finish;
    csv_file_dump fifo_csv_dumper_1019;
    csv_file_dump cstatus_csv_dumper_1019;
    df_fifo_monitor fifo_monitor_1019;
    df_fifo_intf fifo_intf_1020(clock,reset);
    assign fifo_intf_1020.rd_en = AESL_inst_myproject.layer2_out_1019_U.if_read & AESL_inst_myproject.layer2_out_1019_U.if_empty_n;
    assign fifo_intf_1020.wr_en = AESL_inst_myproject.layer2_out_1019_U.if_write & AESL_inst_myproject.layer2_out_1019_U.if_full_n;
    assign fifo_intf_1020.fifo_rd_block = 0;
    assign fifo_intf_1020.fifo_wr_block = 0;
    assign fifo_intf_1020.finish = finish;
    csv_file_dump fifo_csv_dumper_1020;
    csv_file_dump cstatus_csv_dumper_1020;
    df_fifo_monitor fifo_monitor_1020;
    df_fifo_intf fifo_intf_1021(clock,reset);
    assign fifo_intf_1021.rd_en = AESL_inst_myproject.layer2_out_1020_U.if_read & AESL_inst_myproject.layer2_out_1020_U.if_empty_n;
    assign fifo_intf_1021.wr_en = AESL_inst_myproject.layer2_out_1020_U.if_write & AESL_inst_myproject.layer2_out_1020_U.if_full_n;
    assign fifo_intf_1021.fifo_rd_block = 0;
    assign fifo_intf_1021.fifo_wr_block = 0;
    assign fifo_intf_1021.finish = finish;
    csv_file_dump fifo_csv_dumper_1021;
    csv_file_dump cstatus_csv_dumper_1021;
    df_fifo_monitor fifo_monitor_1021;
    df_fifo_intf fifo_intf_1022(clock,reset);
    assign fifo_intf_1022.rd_en = AESL_inst_myproject.layer2_out_1021_U.if_read & AESL_inst_myproject.layer2_out_1021_U.if_empty_n;
    assign fifo_intf_1022.wr_en = AESL_inst_myproject.layer2_out_1021_U.if_write & AESL_inst_myproject.layer2_out_1021_U.if_full_n;
    assign fifo_intf_1022.fifo_rd_block = 0;
    assign fifo_intf_1022.fifo_wr_block = 0;
    assign fifo_intf_1022.finish = finish;
    csv_file_dump fifo_csv_dumper_1022;
    csv_file_dump cstatus_csv_dumper_1022;
    df_fifo_monitor fifo_monitor_1022;
    df_fifo_intf fifo_intf_1023(clock,reset);
    assign fifo_intf_1023.rd_en = AESL_inst_myproject.layer2_out_1022_U.if_read & AESL_inst_myproject.layer2_out_1022_U.if_empty_n;
    assign fifo_intf_1023.wr_en = AESL_inst_myproject.layer2_out_1022_U.if_write & AESL_inst_myproject.layer2_out_1022_U.if_full_n;
    assign fifo_intf_1023.fifo_rd_block = 0;
    assign fifo_intf_1023.fifo_wr_block = 0;
    assign fifo_intf_1023.finish = finish;
    csv_file_dump fifo_csv_dumper_1023;
    csv_file_dump cstatus_csv_dumper_1023;
    df_fifo_monitor fifo_monitor_1023;
    df_fifo_intf fifo_intf_1024(clock,reset);
    assign fifo_intf_1024.rd_en = AESL_inst_myproject.layer2_out_1023_U.if_read & AESL_inst_myproject.layer2_out_1023_U.if_empty_n;
    assign fifo_intf_1024.wr_en = AESL_inst_myproject.layer2_out_1023_U.if_write & AESL_inst_myproject.layer2_out_1023_U.if_full_n;
    assign fifo_intf_1024.fifo_rd_block = 0;
    assign fifo_intf_1024.fifo_wr_block = 0;
    assign fifo_intf_1024.finish = finish;
    csv_file_dump fifo_csv_dumper_1024;
    csv_file_dump cstatus_csv_dumper_1024;
    df_fifo_monitor fifo_monitor_1024;
    df_fifo_intf fifo_intf_1025(clock,reset);
    assign fifo_intf_1025.rd_en = AESL_inst_myproject.layer2_out_1024_U.if_read & AESL_inst_myproject.layer2_out_1024_U.if_empty_n;
    assign fifo_intf_1025.wr_en = AESL_inst_myproject.layer2_out_1024_U.if_write & AESL_inst_myproject.layer2_out_1024_U.if_full_n;
    assign fifo_intf_1025.fifo_rd_block = 0;
    assign fifo_intf_1025.fifo_wr_block = 0;
    assign fifo_intf_1025.finish = finish;
    csv_file_dump fifo_csv_dumper_1025;
    csv_file_dump cstatus_csv_dumper_1025;
    df_fifo_monitor fifo_monitor_1025;
    df_fifo_intf fifo_intf_1026(clock,reset);
    assign fifo_intf_1026.rd_en = AESL_inst_myproject.layer2_out_1025_U.if_read & AESL_inst_myproject.layer2_out_1025_U.if_empty_n;
    assign fifo_intf_1026.wr_en = AESL_inst_myproject.layer2_out_1025_U.if_write & AESL_inst_myproject.layer2_out_1025_U.if_full_n;
    assign fifo_intf_1026.fifo_rd_block = 0;
    assign fifo_intf_1026.fifo_wr_block = 0;
    assign fifo_intf_1026.finish = finish;
    csv_file_dump fifo_csv_dumper_1026;
    csv_file_dump cstatus_csv_dumper_1026;
    df_fifo_monitor fifo_monitor_1026;
    df_fifo_intf fifo_intf_1027(clock,reset);
    assign fifo_intf_1027.rd_en = AESL_inst_myproject.layer2_out_1026_U.if_read & AESL_inst_myproject.layer2_out_1026_U.if_empty_n;
    assign fifo_intf_1027.wr_en = AESL_inst_myproject.layer2_out_1026_U.if_write & AESL_inst_myproject.layer2_out_1026_U.if_full_n;
    assign fifo_intf_1027.fifo_rd_block = 0;
    assign fifo_intf_1027.fifo_wr_block = 0;
    assign fifo_intf_1027.finish = finish;
    csv_file_dump fifo_csv_dumper_1027;
    csv_file_dump cstatus_csv_dumper_1027;
    df_fifo_monitor fifo_monitor_1027;
    df_fifo_intf fifo_intf_1028(clock,reset);
    assign fifo_intf_1028.rd_en = AESL_inst_myproject.layer2_out_1027_U.if_read & AESL_inst_myproject.layer2_out_1027_U.if_empty_n;
    assign fifo_intf_1028.wr_en = AESL_inst_myproject.layer2_out_1027_U.if_write & AESL_inst_myproject.layer2_out_1027_U.if_full_n;
    assign fifo_intf_1028.fifo_rd_block = 0;
    assign fifo_intf_1028.fifo_wr_block = 0;
    assign fifo_intf_1028.finish = finish;
    csv_file_dump fifo_csv_dumper_1028;
    csv_file_dump cstatus_csv_dumper_1028;
    df_fifo_monitor fifo_monitor_1028;
    df_fifo_intf fifo_intf_1029(clock,reset);
    assign fifo_intf_1029.rd_en = AESL_inst_myproject.layer2_out_1028_U.if_read & AESL_inst_myproject.layer2_out_1028_U.if_empty_n;
    assign fifo_intf_1029.wr_en = AESL_inst_myproject.layer2_out_1028_U.if_write & AESL_inst_myproject.layer2_out_1028_U.if_full_n;
    assign fifo_intf_1029.fifo_rd_block = 0;
    assign fifo_intf_1029.fifo_wr_block = 0;
    assign fifo_intf_1029.finish = finish;
    csv_file_dump fifo_csv_dumper_1029;
    csv_file_dump cstatus_csv_dumper_1029;
    df_fifo_monitor fifo_monitor_1029;
    df_fifo_intf fifo_intf_1030(clock,reset);
    assign fifo_intf_1030.rd_en = AESL_inst_myproject.layer2_out_1029_U.if_read & AESL_inst_myproject.layer2_out_1029_U.if_empty_n;
    assign fifo_intf_1030.wr_en = AESL_inst_myproject.layer2_out_1029_U.if_write & AESL_inst_myproject.layer2_out_1029_U.if_full_n;
    assign fifo_intf_1030.fifo_rd_block = 0;
    assign fifo_intf_1030.fifo_wr_block = 0;
    assign fifo_intf_1030.finish = finish;
    csv_file_dump fifo_csv_dumper_1030;
    csv_file_dump cstatus_csv_dumper_1030;
    df_fifo_monitor fifo_monitor_1030;
    df_fifo_intf fifo_intf_1031(clock,reset);
    assign fifo_intf_1031.rd_en = AESL_inst_myproject.layer2_out_1030_U.if_read & AESL_inst_myproject.layer2_out_1030_U.if_empty_n;
    assign fifo_intf_1031.wr_en = AESL_inst_myproject.layer2_out_1030_U.if_write & AESL_inst_myproject.layer2_out_1030_U.if_full_n;
    assign fifo_intf_1031.fifo_rd_block = 0;
    assign fifo_intf_1031.fifo_wr_block = 0;
    assign fifo_intf_1031.finish = finish;
    csv_file_dump fifo_csv_dumper_1031;
    csv_file_dump cstatus_csv_dumper_1031;
    df_fifo_monitor fifo_monitor_1031;
    df_fifo_intf fifo_intf_1032(clock,reset);
    assign fifo_intf_1032.rd_en = AESL_inst_myproject.layer2_out_1031_U.if_read & AESL_inst_myproject.layer2_out_1031_U.if_empty_n;
    assign fifo_intf_1032.wr_en = AESL_inst_myproject.layer2_out_1031_U.if_write & AESL_inst_myproject.layer2_out_1031_U.if_full_n;
    assign fifo_intf_1032.fifo_rd_block = 0;
    assign fifo_intf_1032.fifo_wr_block = 0;
    assign fifo_intf_1032.finish = finish;
    csv_file_dump fifo_csv_dumper_1032;
    csv_file_dump cstatus_csv_dumper_1032;
    df_fifo_monitor fifo_monitor_1032;
    df_fifo_intf fifo_intf_1033(clock,reset);
    assign fifo_intf_1033.rd_en = AESL_inst_myproject.layer2_out_1032_U.if_read & AESL_inst_myproject.layer2_out_1032_U.if_empty_n;
    assign fifo_intf_1033.wr_en = AESL_inst_myproject.layer2_out_1032_U.if_write & AESL_inst_myproject.layer2_out_1032_U.if_full_n;
    assign fifo_intf_1033.fifo_rd_block = 0;
    assign fifo_intf_1033.fifo_wr_block = 0;
    assign fifo_intf_1033.finish = finish;
    csv_file_dump fifo_csv_dumper_1033;
    csv_file_dump cstatus_csv_dumper_1033;
    df_fifo_monitor fifo_monitor_1033;
    df_fifo_intf fifo_intf_1034(clock,reset);
    assign fifo_intf_1034.rd_en = AESL_inst_myproject.layer2_out_1033_U.if_read & AESL_inst_myproject.layer2_out_1033_U.if_empty_n;
    assign fifo_intf_1034.wr_en = AESL_inst_myproject.layer2_out_1033_U.if_write & AESL_inst_myproject.layer2_out_1033_U.if_full_n;
    assign fifo_intf_1034.fifo_rd_block = 0;
    assign fifo_intf_1034.fifo_wr_block = 0;
    assign fifo_intf_1034.finish = finish;
    csv_file_dump fifo_csv_dumper_1034;
    csv_file_dump cstatus_csv_dumper_1034;
    df_fifo_monitor fifo_monitor_1034;
    df_fifo_intf fifo_intf_1035(clock,reset);
    assign fifo_intf_1035.rd_en = AESL_inst_myproject.layer2_out_1034_U.if_read & AESL_inst_myproject.layer2_out_1034_U.if_empty_n;
    assign fifo_intf_1035.wr_en = AESL_inst_myproject.layer2_out_1034_U.if_write & AESL_inst_myproject.layer2_out_1034_U.if_full_n;
    assign fifo_intf_1035.fifo_rd_block = 0;
    assign fifo_intf_1035.fifo_wr_block = 0;
    assign fifo_intf_1035.finish = finish;
    csv_file_dump fifo_csv_dumper_1035;
    csv_file_dump cstatus_csv_dumper_1035;
    df_fifo_monitor fifo_monitor_1035;
    df_fifo_intf fifo_intf_1036(clock,reset);
    assign fifo_intf_1036.rd_en = AESL_inst_myproject.layer2_out_1035_U.if_read & AESL_inst_myproject.layer2_out_1035_U.if_empty_n;
    assign fifo_intf_1036.wr_en = AESL_inst_myproject.layer2_out_1035_U.if_write & AESL_inst_myproject.layer2_out_1035_U.if_full_n;
    assign fifo_intf_1036.fifo_rd_block = 0;
    assign fifo_intf_1036.fifo_wr_block = 0;
    assign fifo_intf_1036.finish = finish;
    csv_file_dump fifo_csv_dumper_1036;
    csv_file_dump cstatus_csv_dumper_1036;
    df_fifo_monitor fifo_monitor_1036;
    df_fifo_intf fifo_intf_1037(clock,reset);
    assign fifo_intf_1037.rd_en = AESL_inst_myproject.layer2_out_1036_U.if_read & AESL_inst_myproject.layer2_out_1036_U.if_empty_n;
    assign fifo_intf_1037.wr_en = AESL_inst_myproject.layer2_out_1036_U.if_write & AESL_inst_myproject.layer2_out_1036_U.if_full_n;
    assign fifo_intf_1037.fifo_rd_block = 0;
    assign fifo_intf_1037.fifo_wr_block = 0;
    assign fifo_intf_1037.finish = finish;
    csv_file_dump fifo_csv_dumper_1037;
    csv_file_dump cstatus_csv_dumper_1037;
    df_fifo_monitor fifo_monitor_1037;
    df_fifo_intf fifo_intf_1038(clock,reset);
    assign fifo_intf_1038.rd_en = AESL_inst_myproject.layer2_out_1037_U.if_read & AESL_inst_myproject.layer2_out_1037_U.if_empty_n;
    assign fifo_intf_1038.wr_en = AESL_inst_myproject.layer2_out_1037_U.if_write & AESL_inst_myproject.layer2_out_1037_U.if_full_n;
    assign fifo_intf_1038.fifo_rd_block = 0;
    assign fifo_intf_1038.fifo_wr_block = 0;
    assign fifo_intf_1038.finish = finish;
    csv_file_dump fifo_csv_dumper_1038;
    csv_file_dump cstatus_csv_dumper_1038;
    df_fifo_monitor fifo_monitor_1038;
    df_fifo_intf fifo_intf_1039(clock,reset);
    assign fifo_intf_1039.rd_en = AESL_inst_myproject.layer2_out_1038_U.if_read & AESL_inst_myproject.layer2_out_1038_U.if_empty_n;
    assign fifo_intf_1039.wr_en = AESL_inst_myproject.layer2_out_1038_U.if_write & AESL_inst_myproject.layer2_out_1038_U.if_full_n;
    assign fifo_intf_1039.fifo_rd_block = 0;
    assign fifo_intf_1039.fifo_wr_block = 0;
    assign fifo_intf_1039.finish = finish;
    csv_file_dump fifo_csv_dumper_1039;
    csv_file_dump cstatus_csv_dumper_1039;
    df_fifo_monitor fifo_monitor_1039;
    df_fifo_intf fifo_intf_1040(clock,reset);
    assign fifo_intf_1040.rd_en = AESL_inst_myproject.layer2_out_1039_U.if_read & AESL_inst_myproject.layer2_out_1039_U.if_empty_n;
    assign fifo_intf_1040.wr_en = AESL_inst_myproject.layer2_out_1039_U.if_write & AESL_inst_myproject.layer2_out_1039_U.if_full_n;
    assign fifo_intf_1040.fifo_rd_block = 0;
    assign fifo_intf_1040.fifo_wr_block = 0;
    assign fifo_intf_1040.finish = finish;
    csv_file_dump fifo_csv_dumper_1040;
    csv_file_dump cstatus_csv_dumper_1040;
    df_fifo_monitor fifo_monitor_1040;
    df_fifo_intf fifo_intf_1041(clock,reset);
    assign fifo_intf_1041.rd_en = AESL_inst_myproject.layer2_out_1040_U.if_read & AESL_inst_myproject.layer2_out_1040_U.if_empty_n;
    assign fifo_intf_1041.wr_en = AESL_inst_myproject.layer2_out_1040_U.if_write & AESL_inst_myproject.layer2_out_1040_U.if_full_n;
    assign fifo_intf_1041.fifo_rd_block = 0;
    assign fifo_intf_1041.fifo_wr_block = 0;
    assign fifo_intf_1041.finish = finish;
    csv_file_dump fifo_csv_dumper_1041;
    csv_file_dump cstatus_csv_dumper_1041;
    df_fifo_monitor fifo_monitor_1041;
    df_fifo_intf fifo_intf_1042(clock,reset);
    assign fifo_intf_1042.rd_en = AESL_inst_myproject.layer2_out_1041_U.if_read & AESL_inst_myproject.layer2_out_1041_U.if_empty_n;
    assign fifo_intf_1042.wr_en = AESL_inst_myproject.layer2_out_1041_U.if_write & AESL_inst_myproject.layer2_out_1041_U.if_full_n;
    assign fifo_intf_1042.fifo_rd_block = 0;
    assign fifo_intf_1042.fifo_wr_block = 0;
    assign fifo_intf_1042.finish = finish;
    csv_file_dump fifo_csv_dumper_1042;
    csv_file_dump cstatus_csv_dumper_1042;
    df_fifo_monitor fifo_monitor_1042;
    df_fifo_intf fifo_intf_1043(clock,reset);
    assign fifo_intf_1043.rd_en = AESL_inst_myproject.layer2_out_1042_U.if_read & AESL_inst_myproject.layer2_out_1042_U.if_empty_n;
    assign fifo_intf_1043.wr_en = AESL_inst_myproject.layer2_out_1042_U.if_write & AESL_inst_myproject.layer2_out_1042_U.if_full_n;
    assign fifo_intf_1043.fifo_rd_block = 0;
    assign fifo_intf_1043.fifo_wr_block = 0;
    assign fifo_intf_1043.finish = finish;
    csv_file_dump fifo_csv_dumper_1043;
    csv_file_dump cstatus_csv_dumper_1043;
    df_fifo_monitor fifo_monitor_1043;
    df_fifo_intf fifo_intf_1044(clock,reset);
    assign fifo_intf_1044.rd_en = AESL_inst_myproject.layer2_out_1043_U.if_read & AESL_inst_myproject.layer2_out_1043_U.if_empty_n;
    assign fifo_intf_1044.wr_en = AESL_inst_myproject.layer2_out_1043_U.if_write & AESL_inst_myproject.layer2_out_1043_U.if_full_n;
    assign fifo_intf_1044.fifo_rd_block = 0;
    assign fifo_intf_1044.fifo_wr_block = 0;
    assign fifo_intf_1044.finish = finish;
    csv_file_dump fifo_csv_dumper_1044;
    csv_file_dump cstatus_csv_dumper_1044;
    df_fifo_monitor fifo_monitor_1044;
    df_fifo_intf fifo_intf_1045(clock,reset);
    assign fifo_intf_1045.rd_en = AESL_inst_myproject.layer2_out_1044_U.if_read & AESL_inst_myproject.layer2_out_1044_U.if_empty_n;
    assign fifo_intf_1045.wr_en = AESL_inst_myproject.layer2_out_1044_U.if_write & AESL_inst_myproject.layer2_out_1044_U.if_full_n;
    assign fifo_intf_1045.fifo_rd_block = 0;
    assign fifo_intf_1045.fifo_wr_block = 0;
    assign fifo_intf_1045.finish = finish;
    csv_file_dump fifo_csv_dumper_1045;
    csv_file_dump cstatus_csv_dumper_1045;
    df_fifo_monitor fifo_monitor_1045;
    df_fifo_intf fifo_intf_1046(clock,reset);
    assign fifo_intf_1046.rd_en = AESL_inst_myproject.layer2_out_1045_U.if_read & AESL_inst_myproject.layer2_out_1045_U.if_empty_n;
    assign fifo_intf_1046.wr_en = AESL_inst_myproject.layer2_out_1045_U.if_write & AESL_inst_myproject.layer2_out_1045_U.if_full_n;
    assign fifo_intf_1046.fifo_rd_block = 0;
    assign fifo_intf_1046.fifo_wr_block = 0;
    assign fifo_intf_1046.finish = finish;
    csv_file_dump fifo_csv_dumper_1046;
    csv_file_dump cstatus_csv_dumper_1046;
    df_fifo_monitor fifo_monitor_1046;
    df_fifo_intf fifo_intf_1047(clock,reset);
    assign fifo_intf_1047.rd_en = AESL_inst_myproject.layer2_out_1046_U.if_read & AESL_inst_myproject.layer2_out_1046_U.if_empty_n;
    assign fifo_intf_1047.wr_en = AESL_inst_myproject.layer2_out_1046_U.if_write & AESL_inst_myproject.layer2_out_1046_U.if_full_n;
    assign fifo_intf_1047.fifo_rd_block = 0;
    assign fifo_intf_1047.fifo_wr_block = 0;
    assign fifo_intf_1047.finish = finish;
    csv_file_dump fifo_csv_dumper_1047;
    csv_file_dump cstatus_csv_dumper_1047;
    df_fifo_monitor fifo_monitor_1047;
    df_fifo_intf fifo_intf_1048(clock,reset);
    assign fifo_intf_1048.rd_en = AESL_inst_myproject.layer2_out_1047_U.if_read & AESL_inst_myproject.layer2_out_1047_U.if_empty_n;
    assign fifo_intf_1048.wr_en = AESL_inst_myproject.layer2_out_1047_U.if_write & AESL_inst_myproject.layer2_out_1047_U.if_full_n;
    assign fifo_intf_1048.fifo_rd_block = 0;
    assign fifo_intf_1048.fifo_wr_block = 0;
    assign fifo_intf_1048.finish = finish;
    csv_file_dump fifo_csv_dumper_1048;
    csv_file_dump cstatus_csv_dumper_1048;
    df_fifo_monitor fifo_monitor_1048;
    df_fifo_intf fifo_intf_1049(clock,reset);
    assign fifo_intf_1049.rd_en = AESL_inst_myproject.layer2_out_1048_U.if_read & AESL_inst_myproject.layer2_out_1048_U.if_empty_n;
    assign fifo_intf_1049.wr_en = AESL_inst_myproject.layer2_out_1048_U.if_write & AESL_inst_myproject.layer2_out_1048_U.if_full_n;
    assign fifo_intf_1049.fifo_rd_block = 0;
    assign fifo_intf_1049.fifo_wr_block = 0;
    assign fifo_intf_1049.finish = finish;
    csv_file_dump fifo_csv_dumper_1049;
    csv_file_dump cstatus_csv_dumper_1049;
    df_fifo_monitor fifo_monitor_1049;
    df_fifo_intf fifo_intf_1050(clock,reset);
    assign fifo_intf_1050.rd_en = AESL_inst_myproject.layer2_out_1049_U.if_read & AESL_inst_myproject.layer2_out_1049_U.if_empty_n;
    assign fifo_intf_1050.wr_en = AESL_inst_myproject.layer2_out_1049_U.if_write & AESL_inst_myproject.layer2_out_1049_U.if_full_n;
    assign fifo_intf_1050.fifo_rd_block = 0;
    assign fifo_intf_1050.fifo_wr_block = 0;
    assign fifo_intf_1050.finish = finish;
    csv_file_dump fifo_csv_dumper_1050;
    csv_file_dump cstatus_csv_dumper_1050;
    df_fifo_monitor fifo_monitor_1050;
    df_fifo_intf fifo_intf_1051(clock,reset);
    assign fifo_intf_1051.rd_en = AESL_inst_myproject.layer2_out_1050_U.if_read & AESL_inst_myproject.layer2_out_1050_U.if_empty_n;
    assign fifo_intf_1051.wr_en = AESL_inst_myproject.layer2_out_1050_U.if_write & AESL_inst_myproject.layer2_out_1050_U.if_full_n;
    assign fifo_intf_1051.fifo_rd_block = 0;
    assign fifo_intf_1051.fifo_wr_block = 0;
    assign fifo_intf_1051.finish = finish;
    csv_file_dump fifo_csv_dumper_1051;
    csv_file_dump cstatus_csv_dumper_1051;
    df_fifo_monitor fifo_monitor_1051;
    df_fifo_intf fifo_intf_1052(clock,reset);
    assign fifo_intf_1052.rd_en = AESL_inst_myproject.layer2_out_1051_U.if_read & AESL_inst_myproject.layer2_out_1051_U.if_empty_n;
    assign fifo_intf_1052.wr_en = AESL_inst_myproject.layer2_out_1051_U.if_write & AESL_inst_myproject.layer2_out_1051_U.if_full_n;
    assign fifo_intf_1052.fifo_rd_block = 0;
    assign fifo_intf_1052.fifo_wr_block = 0;
    assign fifo_intf_1052.finish = finish;
    csv_file_dump fifo_csv_dumper_1052;
    csv_file_dump cstatus_csv_dumper_1052;
    df_fifo_monitor fifo_monitor_1052;
    df_fifo_intf fifo_intf_1053(clock,reset);
    assign fifo_intf_1053.rd_en = AESL_inst_myproject.layer2_out_1052_U.if_read & AESL_inst_myproject.layer2_out_1052_U.if_empty_n;
    assign fifo_intf_1053.wr_en = AESL_inst_myproject.layer2_out_1052_U.if_write & AESL_inst_myproject.layer2_out_1052_U.if_full_n;
    assign fifo_intf_1053.fifo_rd_block = 0;
    assign fifo_intf_1053.fifo_wr_block = 0;
    assign fifo_intf_1053.finish = finish;
    csv_file_dump fifo_csv_dumper_1053;
    csv_file_dump cstatus_csv_dumper_1053;
    df_fifo_monitor fifo_monitor_1053;
    df_fifo_intf fifo_intf_1054(clock,reset);
    assign fifo_intf_1054.rd_en = AESL_inst_myproject.layer2_out_1053_U.if_read & AESL_inst_myproject.layer2_out_1053_U.if_empty_n;
    assign fifo_intf_1054.wr_en = AESL_inst_myproject.layer2_out_1053_U.if_write & AESL_inst_myproject.layer2_out_1053_U.if_full_n;
    assign fifo_intf_1054.fifo_rd_block = 0;
    assign fifo_intf_1054.fifo_wr_block = 0;
    assign fifo_intf_1054.finish = finish;
    csv_file_dump fifo_csv_dumper_1054;
    csv_file_dump cstatus_csv_dumper_1054;
    df_fifo_monitor fifo_monitor_1054;
    df_fifo_intf fifo_intf_1055(clock,reset);
    assign fifo_intf_1055.rd_en = AESL_inst_myproject.layer2_out_1054_U.if_read & AESL_inst_myproject.layer2_out_1054_U.if_empty_n;
    assign fifo_intf_1055.wr_en = AESL_inst_myproject.layer2_out_1054_U.if_write & AESL_inst_myproject.layer2_out_1054_U.if_full_n;
    assign fifo_intf_1055.fifo_rd_block = 0;
    assign fifo_intf_1055.fifo_wr_block = 0;
    assign fifo_intf_1055.finish = finish;
    csv_file_dump fifo_csv_dumper_1055;
    csv_file_dump cstatus_csv_dumper_1055;
    df_fifo_monitor fifo_monitor_1055;
    df_fifo_intf fifo_intf_1056(clock,reset);
    assign fifo_intf_1056.rd_en = AESL_inst_myproject.layer2_out_1055_U.if_read & AESL_inst_myproject.layer2_out_1055_U.if_empty_n;
    assign fifo_intf_1056.wr_en = AESL_inst_myproject.layer2_out_1055_U.if_write & AESL_inst_myproject.layer2_out_1055_U.if_full_n;
    assign fifo_intf_1056.fifo_rd_block = 0;
    assign fifo_intf_1056.fifo_wr_block = 0;
    assign fifo_intf_1056.finish = finish;
    csv_file_dump fifo_csv_dumper_1056;
    csv_file_dump cstatus_csv_dumper_1056;
    df_fifo_monitor fifo_monitor_1056;
    df_fifo_intf fifo_intf_1057(clock,reset);
    assign fifo_intf_1057.rd_en = AESL_inst_myproject.layer2_out_1056_U.if_read & AESL_inst_myproject.layer2_out_1056_U.if_empty_n;
    assign fifo_intf_1057.wr_en = AESL_inst_myproject.layer2_out_1056_U.if_write & AESL_inst_myproject.layer2_out_1056_U.if_full_n;
    assign fifo_intf_1057.fifo_rd_block = 0;
    assign fifo_intf_1057.fifo_wr_block = 0;
    assign fifo_intf_1057.finish = finish;
    csv_file_dump fifo_csv_dumper_1057;
    csv_file_dump cstatus_csv_dumper_1057;
    df_fifo_monitor fifo_monitor_1057;
    df_fifo_intf fifo_intf_1058(clock,reset);
    assign fifo_intf_1058.rd_en = AESL_inst_myproject.layer2_out_1057_U.if_read & AESL_inst_myproject.layer2_out_1057_U.if_empty_n;
    assign fifo_intf_1058.wr_en = AESL_inst_myproject.layer2_out_1057_U.if_write & AESL_inst_myproject.layer2_out_1057_U.if_full_n;
    assign fifo_intf_1058.fifo_rd_block = 0;
    assign fifo_intf_1058.fifo_wr_block = 0;
    assign fifo_intf_1058.finish = finish;
    csv_file_dump fifo_csv_dumper_1058;
    csv_file_dump cstatus_csv_dumper_1058;
    df_fifo_monitor fifo_monitor_1058;
    df_fifo_intf fifo_intf_1059(clock,reset);
    assign fifo_intf_1059.rd_en = AESL_inst_myproject.layer2_out_1058_U.if_read & AESL_inst_myproject.layer2_out_1058_U.if_empty_n;
    assign fifo_intf_1059.wr_en = AESL_inst_myproject.layer2_out_1058_U.if_write & AESL_inst_myproject.layer2_out_1058_U.if_full_n;
    assign fifo_intf_1059.fifo_rd_block = 0;
    assign fifo_intf_1059.fifo_wr_block = 0;
    assign fifo_intf_1059.finish = finish;
    csv_file_dump fifo_csv_dumper_1059;
    csv_file_dump cstatus_csv_dumper_1059;
    df_fifo_monitor fifo_monitor_1059;
    df_fifo_intf fifo_intf_1060(clock,reset);
    assign fifo_intf_1060.rd_en = AESL_inst_myproject.layer2_out_1059_U.if_read & AESL_inst_myproject.layer2_out_1059_U.if_empty_n;
    assign fifo_intf_1060.wr_en = AESL_inst_myproject.layer2_out_1059_U.if_write & AESL_inst_myproject.layer2_out_1059_U.if_full_n;
    assign fifo_intf_1060.fifo_rd_block = 0;
    assign fifo_intf_1060.fifo_wr_block = 0;
    assign fifo_intf_1060.finish = finish;
    csv_file_dump fifo_csv_dumper_1060;
    csv_file_dump cstatus_csv_dumper_1060;
    df_fifo_monitor fifo_monitor_1060;
    df_fifo_intf fifo_intf_1061(clock,reset);
    assign fifo_intf_1061.rd_en = AESL_inst_myproject.layer2_out_1060_U.if_read & AESL_inst_myproject.layer2_out_1060_U.if_empty_n;
    assign fifo_intf_1061.wr_en = AESL_inst_myproject.layer2_out_1060_U.if_write & AESL_inst_myproject.layer2_out_1060_U.if_full_n;
    assign fifo_intf_1061.fifo_rd_block = 0;
    assign fifo_intf_1061.fifo_wr_block = 0;
    assign fifo_intf_1061.finish = finish;
    csv_file_dump fifo_csv_dumper_1061;
    csv_file_dump cstatus_csv_dumper_1061;
    df_fifo_monitor fifo_monitor_1061;
    df_fifo_intf fifo_intf_1062(clock,reset);
    assign fifo_intf_1062.rd_en = AESL_inst_myproject.layer2_out_1061_U.if_read & AESL_inst_myproject.layer2_out_1061_U.if_empty_n;
    assign fifo_intf_1062.wr_en = AESL_inst_myproject.layer2_out_1061_U.if_write & AESL_inst_myproject.layer2_out_1061_U.if_full_n;
    assign fifo_intf_1062.fifo_rd_block = 0;
    assign fifo_intf_1062.fifo_wr_block = 0;
    assign fifo_intf_1062.finish = finish;
    csv_file_dump fifo_csv_dumper_1062;
    csv_file_dump cstatus_csv_dumper_1062;
    df_fifo_monitor fifo_monitor_1062;
    df_fifo_intf fifo_intf_1063(clock,reset);
    assign fifo_intf_1063.rd_en = AESL_inst_myproject.layer2_out_1062_U.if_read & AESL_inst_myproject.layer2_out_1062_U.if_empty_n;
    assign fifo_intf_1063.wr_en = AESL_inst_myproject.layer2_out_1062_U.if_write & AESL_inst_myproject.layer2_out_1062_U.if_full_n;
    assign fifo_intf_1063.fifo_rd_block = 0;
    assign fifo_intf_1063.fifo_wr_block = 0;
    assign fifo_intf_1063.finish = finish;
    csv_file_dump fifo_csv_dumper_1063;
    csv_file_dump cstatus_csv_dumper_1063;
    df_fifo_monitor fifo_monitor_1063;
    df_fifo_intf fifo_intf_1064(clock,reset);
    assign fifo_intf_1064.rd_en = AESL_inst_myproject.layer2_out_1063_U.if_read & AESL_inst_myproject.layer2_out_1063_U.if_empty_n;
    assign fifo_intf_1064.wr_en = AESL_inst_myproject.layer2_out_1063_U.if_write & AESL_inst_myproject.layer2_out_1063_U.if_full_n;
    assign fifo_intf_1064.fifo_rd_block = 0;
    assign fifo_intf_1064.fifo_wr_block = 0;
    assign fifo_intf_1064.finish = finish;
    csv_file_dump fifo_csv_dumper_1064;
    csv_file_dump cstatus_csv_dumper_1064;
    df_fifo_monitor fifo_monitor_1064;
    df_fifo_intf fifo_intf_1065(clock,reset);
    assign fifo_intf_1065.rd_en = AESL_inst_myproject.layer2_out_1064_U.if_read & AESL_inst_myproject.layer2_out_1064_U.if_empty_n;
    assign fifo_intf_1065.wr_en = AESL_inst_myproject.layer2_out_1064_U.if_write & AESL_inst_myproject.layer2_out_1064_U.if_full_n;
    assign fifo_intf_1065.fifo_rd_block = 0;
    assign fifo_intf_1065.fifo_wr_block = 0;
    assign fifo_intf_1065.finish = finish;
    csv_file_dump fifo_csv_dumper_1065;
    csv_file_dump cstatus_csv_dumper_1065;
    df_fifo_monitor fifo_monitor_1065;
    df_fifo_intf fifo_intf_1066(clock,reset);
    assign fifo_intf_1066.rd_en = AESL_inst_myproject.layer2_out_1065_U.if_read & AESL_inst_myproject.layer2_out_1065_U.if_empty_n;
    assign fifo_intf_1066.wr_en = AESL_inst_myproject.layer2_out_1065_U.if_write & AESL_inst_myproject.layer2_out_1065_U.if_full_n;
    assign fifo_intf_1066.fifo_rd_block = 0;
    assign fifo_intf_1066.fifo_wr_block = 0;
    assign fifo_intf_1066.finish = finish;
    csv_file_dump fifo_csv_dumper_1066;
    csv_file_dump cstatus_csv_dumper_1066;
    df_fifo_monitor fifo_monitor_1066;
    df_fifo_intf fifo_intf_1067(clock,reset);
    assign fifo_intf_1067.rd_en = AESL_inst_myproject.layer2_out_1066_U.if_read & AESL_inst_myproject.layer2_out_1066_U.if_empty_n;
    assign fifo_intf_1067.wr_en = AESL_inst_myproject.layer2_out_1066_U.if_write & AESL_inst_myproject.layer2_out_1066_U.if_full_n;
    assign fifo_intf_1067.fifo_rd_block = 0;
    assign fifo_intf_1067.fifo_wr_block = 0;
    assign fifo_intf_1067.finish = finish;
    csv_file_dump fifo_csv_dumper_1067;
    csv_file_dump cstatus_csv_dumper_1067;
    df_fifo_monitor fifo_monitor_1067;
    df_fifo_intf fifo_intf_1068(clock,reset);
    assign fifo_intf_1068.rd_en = AESL_inst_myproject.layer2_out_1067_U.if_read & AESL_inst_myproject.layer2_out_1067_U.if_empty_n;
    assign fifo_intf_1068.wr_en = AESL_inst_myproject.layer2_out_1067_U.if_write & AESL_inst_myproject.layer2_out_1067_U.if_full_n;
    assign fifo_intf_1068.fifo_rd_block = 0;
    assign fifo_intf_1068.fifo_wr_block = 0;
    assign fifo_intf_1068.finish = finish;
    csv_file_dump fifo_csv_dumper_1068;
    csv_file_dump cstatus_csv_dumper_1068;
    df_fifo_monitor fifo_monitor_1068;
    df_fifo_intf fifo_intf_1069(clock,reset);
    assign fifo_intf_1069.rd_en = AESL_inst_myproject.layer2_out_1068_U.if_read & AESL_inst_myproject.layer2_out_1068_U.if_empty_n;
    assign fifo_intf_1069.wr_en = AESL_inst_myproject.layer2_out_1068_U.if_write & AESL_inst_myproject.layer2_out_1068_U.if_full_n;
    assign fifo_intf_1069.fifo_rd_block = 0;
    assign fifo_intf_1069.fifo_wr_block = 0;
    assign fifo_intf_1069.finish = finish;
    csv_file_dump fifo_csv_dumper_1069;
    csv_file_dump cstatus_csv_dumper_1069;
    df_fifo_monitor fifo_monitor_1069;
    df_fifo_intf fifo_intf_1070(clock,reset);
    assign fifo_intf_1070.rd_en = AESL_inst_myproject.layer2_out_1069_U.if_read & AESL_inst_myproject.layer2_out_1069_U.if_empty_n;
    assign fifo_intf_1070.wr_en = AESL_inst_myproject.layer2_out_1069_U.if_write & AESL_inst_myproject.layer2_out_1069_U.if_full_n;
    assign fifo_intf_1070.fifo_rd_block = 0;
    assign fifo_intf_1070.fifo_wr_block = 0;
    assign fifo_intf_1070.finish = finish;
    csv_file_dump fifo_csv_dumper_1070;
    csv_file_dump cstatus_csv_dumper_1070;
    df_fifo_monitor fifo_monitor_1070;
    df_fifo_intf fifo_intf_1071(clock,reset);
    assign fifo_intf_1071.rd_en = AESL_inst_myproject.layer2_out_1070_U.if_read & AESL_inst_myproject.layer2_out_1070_U.if_empty_n;
    assign fifo_intf_1071.wr_en = AESL_inst_myproject.layer2_out_1070_U.if_write & AESL_inst_myproject.layer2_out_1070_U.if_full_n;
    assign fifo_intf_1071.fifo_rd_block = 0;
    assign fifo_intf_1071.fifo_wr_block = 0;
    assign fifo_intf_1071.finish = finish;
    csv_file_dump fifo_csv_dumper_1071;
    csv_file_dump cstatus_csv_dumper_1071;
    df_fifo_monitor fifo_monitor_1071;
    df_fifo_intf fifo_intf_1072(clock,reset);
    assign fifo_intf_1072.rd_en = AESL_inst_myproject.layer2_out_1071_U.if_read & AESL_inst_myproject.layer2_out_1071_U.if_empty_n;
    assign fifo_intf_1072.wr_en = AESL_inst_myproject.layer2_out_1071_U.if_write & AESL_inst_myproject.layer2_out_1071_U.if_full_n;
    assign fifo_intf_1072.fifo_rd_block = 0;
    assign fifo_intf_1072.fifo_wr_block = 0;
    assign fifo_intf_1072.finish = finish;
    csv_file_dump fifo_csv_dumper_1072;
    csv_file_dump cstatus_csv_dumper_1072;
    df_fifo_monitor fifo_monitor_1072;
    df_fifo_intf fifo_intf_1073(clock,reset);
    assign fifo_intf_1073.rd_en = AESL_inst_myproject.layer2_out_1072_U.if_read & AESL_inst_myproject.layer2_out_1072_U.if_empty_n;
    assign fifo_intf_1073.wr_en = AESL_inst_myproject.layer2_out_1072_U.if_write & AESL_inst_myproject.layer2_out_1072_U.if_full_n;
    assign fifo_intf_1073.fifo_rd_block = 0;
    assign fifo_intf_1073.fifo_wr_block = 0;
    assign fifo_intf_1073.finish = finish;
    csv_file_dump fifo_csv_dumper_1073;
    csv_file_dump cstatus_csv_dumper_1073;
    df_fifo_monitor fifo_monitor_1073;
    df_fifo_intf fifo_intf_1074(clock,reset);
    assign fifo_intf_1074.rd_en = AESL_inst_myproject.layer2_out_1073_U.if_read & AESL_inst_myproject.layer2_out_1073_U.if_empty_n;
    assign fifo_intf_1074.wr_en = AESL_inst_myproject.layer2_out_1073_U.if_write & AESL_inst_myproject.layer2_out_1073_U.if_full_n;
    assign fifo_intf_1074.fifo_rd_block = 0;
    assign fifo_intf_1074.fifo_wr_block = 0;
    assign fifo_intf_1074.finish = finish;
    csv_file_dump fifo_csv_dumper_1074;
    csv_file_dump cstatus_csv_dumper_1074;
    df_fifo_monitor fifo_monitor_1074;
    df_fifo_intf fifo_intf_1075(clock,reset);
    assign fifo_intf_1075.rd_en = AESL_inst_myproject.layer2_out_1074_U.if_read & AESL_inst_myproject.layer2_out_1074_U.if_empty_n;
    assign fifo_intf_1075.wr_en = AESL_inst_myproject.layer2_out_1074_U.if_write & AESL_inst_myproject.layer2_out_1074_U.if_full_n;
    assign fifo_intf_1075.fifo_rd_block = 0;
    assign fifo_intf_1075.fifo_wr_block = 0;
    assign fifo_intf_1075.finish = finish;
    csv_file_dump fifo_csv_dumper_1075;
    csv_file_dump cstatus_csv_dumper_1075;
    df_fifo_monitor fifo_monitor_1075;
    df_fifo_intf fifo_intf_1076(clock,reset);
    assign fifo_intf_1076.rd_en = AESL_inst_myproject.layer2_out_1075_U.if_read & AESL_inst_myproject.layer2_out_1075_U.if_empty_n;
    assign fifo_intf_1076.wr_en = AESL_inst_myproject.layer2_out_1075_U.if_write & AESL_inst_myproject.layer2_out_1075_U.if_full_n;
    assign fifo_intf_1076.fifo_rd_block = 0;
    assign fifo_intf_1076.fifo_wr_block = 0;
    assign fifo_intf_1076.finish = finish;
    csv_file_dump fifo_csv_dumper_1076;
    csv_file_dump cstatus_csv_dumper_1076;
    df_fifo_monitor fifo_monitor_1076;
    df_fifo_intf fifo_intf_1077(clock,reset);
    assign fifo_intf_1077.rd_en = AESL_inst_myproject.layer2_out_1076_U.if_read & AESL_inst_myproject.layer2_out_1076_U.if_empty_n;
    assign fifo_intf_1077.wr_en = AESL_inst_myproject.layer2_out_1076_U.if_write & AESL_inst_myproject.layer2_out_1076_U.if_full_n;
    assign fifo_intf_1077.fifo_rd_block = 0;
    assign fifo_intf_1077.fifo_wr_block = 0;
    assign fifo_intf_1077.finish = finish;
    csv_file_dump fifo_csv_dumper_1077;
    csv_file_dump cstatus_csv_dumper_1077;
    df_fifo_monitor fifo_monitor_1077;
    df_fifo_intf fifo_intf_1078(clock,reset);
    assign fifo_intf_1078.rd_en = AESL_inst_myproject.layer2_out_1077_U.if_read & AESL_inst_myproject.layer2_out_1077_U.if_empty_n;
    assign fifo_intf_1078.wr_en = AESL_inst_myproject.layer2_out_1077_U.if_write & AESL_inst_myproject.layer2_out_1077_U.if_full_n;
    assign fifo_intf_1078.fifo_rd_block = 0;
    assign fifo_intf_1078.fifo_wr_block = 0;
    assign fifo_intf_1078.finish = finish;
    csv_file_dump fifo_csv_dumper_1078;
    csv_file_dump cstatus_csv_dumper_1078;
    df_fifo_monitor fifo_monitor_1078;
    df_fifo_intf fifo_intf_1079(clock,reset);
    assign fifo_intf_1079.rd_en = AESL_inst_myproject.layer2_out_1078_U.if_read & AESL_inst_myproject.layer2_out_1078_U.if_empty_n;
    assign fifo_intf_1079.wr_en = AESL_inst_myproject.layer2_out_1078_U.if_write & AESL_inst_myproject.layer2_out_1078_U.if_full_n;
    assign fifo_intf_1079.fifo_rd_block = 0;
    assign fifo_intf_1079.fifo_wr_block = 0;
    assign fifo_intf_1079.finish = finish;
    csv_file_dump fifo_csv_dumper_1079;
    csv_file_dump cstatus_csv_dumper_1079;
    df_fifo_monitor fifo_monitor_1079;
    df_fifo_intf fifo_intf_1080(clock,reset);
    assign fifo_intf_1080.rd_en = AESL_inst_myproject.layer2_out_1079_U.if_read & AESL_inst_myproject.layer2_out_1079_U.if_empty_n;
    assign fifo_intf_1080.wr_en = AESL_inst_myproject.layer2_out_1079_U.if_write & AESL_inst_myproject.layer2_out_1079_U.if_full_n;
    assign fifo_intf_1080.fifo_rd_block = 0;
    assign fifo_intf_1080.fifo_wr_block = 0;
    assign fifo_intf_1080.finish = finish;
    csv_file_dump fifo_csv_dumper_1080;
    csv_file_dump cstatus_csv_dumper_1080;
    df_fifo_monitor fifo_monitor_1080;
    df_fifo_intf fifo_intf_1081(clock,reset);
    assign fifo_intf_1081.rd_en = AESL_inst_myproject.layer2_out_1080_U.if_read & AESL_inst_myproject.layer2_out_1080_U.if_empty_n;
    assign fifo_intf_1081.wr_en = AESL_inst_myproject.layer2_out_1080_U.if_write & AESL_inst_myproject.layer2_out_1080_U.if_full_n;
    assign fifo_intf_1081.fifo_rd_block = 0;
    assign fifo_intf_1081.fifo_wr_block = 0;
    assign fifo_intf_1081.finish = finish;
    csv_file_dump fifo_csv_dumper_1081;
    csv_file_dump cstatus_csv_dumper_1081;
    df_fifo_monitor fifo_monitor_1081;
    df_fifo_intf fifo_intf_1082(clock,reset);
    assign fifo_intf_1082.rd_en = AESL_inst_myproject.layer2_out_1081_U.if_read & AESL_inst_myproject.layer2_out_1081_U.if_empty_n;
    assign fifo_intf_1082.wr_en = AESL_inst_myproject.layer2_out_1081_U.if_write & AESL_inst_myproject.layer2_out_1081_U.if_full_n;
    assign fifo_intf_1082.fifo_rd_block = 0;
    assign fifo_intf_1082.fifo_wr_block = 0;
    assign fifo_intf_1082.finish = finish;
    csv_file_dump fifo_csv_dumper_1082;
    csv_file_dump cstatus_csv_dumper_1082;
    df_fifo_monitor fifo_monitor_1082;
    df_fifo_intf fifo_intf_1083(clock,reset);
    assign fifo_intf_1083.rd_en = AESL_inst_myproject.layer2_out_1082_U.if_read & AESL_inst_myproject.layer2_out_1082_U.if_empty_n;
    assign fifo_intf_1083.wr_en = AESL_inst_myproject.layer2_out_1082_U.if_write & AESL_inst_myproject.layer2_out_1082_U.if_full_n;
    assign fifo_intf_1083.fifo_rd_block = 0;
    assign fifo_intf_1083.fifo_wr_block = 0;
    assign fifo_intf_1083.finish = finish;
    csv_file_dump fifo_csv_dumper_1083;
    csv_file_dump cstatus_csv_dumper_1083;
    df_fifo_monitor fifo_monitor_1083;
    df_fifo_intf fifo_intf_1084(clock,reset);
    assign fifo_intf_1084.rd_en = AESL_inst_myproject.layer2_out_1083_U.if_read & AESL_inst_myproject.layer2_out_1083_U.if_empty_n;
    assign fifo_intf_1084.wr_en = AESL_inst_myproject.layer2_out_1083_U.if_write & AESL_inst_myproject.layer2_out_1083_U.if_full_n;
    assign fifo_intf_1084.fifo_rd_block = 0;
    assign fifo_intf_1084.fifo_wr_block = 0;
    assign fifo_intf_1084.finish = finish;
    csv_file_dump fifo_csv_dumper_1084;
    csv_file_dump cstatus_csv_dumper_1084;
    df_fifo_monitor fifo_monitor_1084;
    df_fifo_intf fifo_intf_1085(clock,reset);
    assign fifo_intf_1085.rd_en = AESL_inst_myproject.layer2_out_1084_U.if_read & AESL_inst_myproject.layer2_out_1084_U.if_empty_n;
    assign fifo_intf_1085.wr_en = AESL_inst_myproject.layer2_out_1084_U.if_write & AESL_inst_myproject.layer2_out_1084_U.if_full_n;
    assign fifo_intf_1085.fifo_rd_block = 0;
    assign fifo_intf_1085.fifo_wr_block = 0;
    assign fifo_intf_1085.finish = finish;
    csv_file_dump fifo_csv_dumper_1085;
    csv_file_dump cstatus_csv_dumper_1085;
    df_fifo_monitor fifo_monitor_1085;
    df_fifo_intf fifo_intf_1086(clock,reset);
    assign fifo_intf_1086.rd_en = AESL_inst_myproject.layer2_out_1085_U.if_read & AESL_inst_myproject.layer2_out_1085_U.if_empty_n;
    assign fifo_intf_1086.wr_en = AESL_inst_myproject.layer2_out_1085_U.if_write & AESL_inst_myproject.layer2_out_1085_U.if_full_n;
    assign fifo_intf_1086.fifo_rd_block = 0;
    assign fifo_intf_1086.fifo_wr_block = 0;
    assign fifo_intf_1086.finish = finish;
    csv_file_dump fifo_csv_dumper_1086;
    csv_file_dump cstatus_csv_dumper_1086;
    df_fifo_monitor fifo_monitor_1086;
    df_fifo_intf fifo_intf_1087(clock,reset);
    assign fifo_intf_1087.rd_en = AESL_inst_myproject.layer2_out_1086_U.if_read & AESL_inst_myproject.layer2_out_1086_U.if_empty_n;
    assign fifo_intf_1087.wr_en = AESL_inst_myproject.layer2_out_1086_U.if_write & AESL_inst_myproject.layer2_out_1086_U.if_full_n;
    assign fifo_intf_1087.fifo_rd_block = 0;
    assign fifo_intf_1087.fifo_wr_block = 0;
    assign fifo_intf_1087.finish = finish;
    csv_file_dump fifo_csv_dumper_1087;
    csv_file_dump cstatus_csv_dumper_1087;
    df_fifo_monitor fifo_monitor_1087;
    df_fifo_intf fifo_intf_1088(clock,reset);
    assign fifo_intf_1088.rd_en = AESL_inst_myproject.layer2_out_1087_U.if_read & AESL_inst_myproject.layer2_out_1087_U.if_empty_n;
    assign fifo_intf_1088.wr_en = AESL_inst_myproject.layer2_out_1087_U.if_write & AESL_inst_myproject.layer2_out_1087_U.if_full_n;
    assign fifo_intf_1088.fifo_rd_block = 0;
    assign fifo_intf_1088.fifo_wr_block = 0;
    assign fifo_intf_1088.finish = finish;
    csv_file_dump fifo_csv_dumper_1088;
    csv_file_dump cstatus_csv_dumper_1088;
    df_fifo_monitor fifo_monitor_1088;
    df_fifo_intf fifo_intf_1089(clock,reset);
    assign fifo_intf_1089.rd_en = AESL_inst_myproject.layer2_out_1088_U.if_read & AESL_inst_myproject.layer2_out_1088_U.if_empty_n;
    assign fifo_intf_1089.wr_en = AESL_inst_myproject.layer2_out_1088_U.if_write & AESL_inst_myproject.layer2_out_1088_U.if_full_n;
    assign fifo_intf_1089.fifo_rd_block = 0;
    assign fifo_intf_1089.fifo_wr_block = 0;
    assign fifo_intf_1089.finish = finish;
    csv_file_dump fifo_csv_dumper_1089;
    csv_file_dump cstatus_csv_dumper_1089;
    df_fifo_monitor fifo_monitor_1089;
    df_fifo_intf fifo_intf_1090(clock,reset);
    assign fifo_intf_1090.rd_en = AESL_inst_myproject.layer2_out_1089_U.if_read & AESL_inst_myproject.layer2_out_1089_U.if_empty_n;
    assign fifo_intf_1090.wr_en = AESL_inst_myproject.layer2_out_1089_U.if_write & AESL_inst_myproject.layer2_out_1089_U.if_full_n;
    assign fifo_intf_1090.fifo_rd_block = 0;
    assign fifo_intf_1090.fifo_wr_block = 0;
    assign fifo_intf_1090.finish = finish;
    csv_file_dump fifo_csv_dumper_1090;
    csv_file_dump cstatus_csv_dumper_1090;
    df_fifo_monitor fifo_monitor_1090;
    df_fifo_intf fifo_intf_1091(clock,reset);
    assign fifo_intf_1091.rd_en = AESL_inst_myproject.layer2_out_1090_U.if_read & AESL_inst_myproject.layer2_out_1090_U.if_empty_n;
    assign fifo_intf_1091.wr_en = AESL_inst_myproject.layer2_out_1090_U.if_write & AESL_inst_myproject.layer2_out_1090_U.if_full_n;
    assign fifo_intf_1091.fifo_rd_block = 0;
    assign fifo_intf_1091.fifo_wr_block = 0;
    assign fifo_intf_1091.finish = finish;
    csv_file_dump fifo_csv_dumper_1091;
    csv_file_dump cstatus_csv_dumper_1091;
    df_fifo_monitor fifo_monitor_1091;
    df_fifo_intf fifo_intf_1092(clock,reset);
    assign fifo_intf_1092.rd_en = AESL_inst_myproject.layer2_out_1091_U.if_read & AESL_inst_myproject.layer2_out_1091_U.if_empty_n;
    assign fifo_intf_1092.wr_en = AESL_inst_myproject.layer2_out_1091_U.if_write & AESL_inst_myproject.layer2_out_1091_U.if_full_n;
    assign fifo_intf_1092.fifo_rd_block = 0;
    assign fifo_intf_1092.fifo_wr_block = 0;
    assign fifo_intf_1092.finish = finish;
    csv_file_dump fifo_csv_dumper_1092;
    csv_file_dump cstatus_csv_dumper_1092;
    df_fifo_monitor fifo_monitor_1092;
    df_fifo_intf fifo_intf_1093(clock,reset);
    assign fifo_intf_1093.rd_en = AESL_inst_myproject.layer2_out_1092_U.if_read & AESL_inst_myproject.layer2_out_1092_U.if_empty_n;
    assign fifo_intf_1093.wr_en = AESL_inst_myproject.layer2_out_1092_U.if_write & AESL_inst_myproject.layer2_out_1092_U.if_full_n;
    assign fifo_intf_1093.fifo_rd_block = 0;
    assign fifo_intf_1093.fifo_wr_block = 0;
    assign fifo_intf_1093.finish = finish;
    csv_file_dump fifo_csv_dumper_1093;
    csv_file_dump cstatus_csv_dumper_1093;
    df_fifo_monitor fifo_monitor_1093;
    df_fifo_intf fifo_intf_1094(clock,reset);
    assign fifo_intf_1094.rd_en = AESL_inst_myproject.layer2_out_1093_U.if_read & AESL_inst_myproject.layer2_out_1093_U.if_empty_n;
    assign fifo_intf_1094.wr_en = AESL_inst_myproject.layer2_out_1093_U.if_write & AESL_inst_myproject.layer2_out_1093_U.if_full_n;
    assign fifo_intf_1094.fifo_rd_block = 0;
    assign fifo_intf_1094.fifo_wr_block = 0;
    assign fifo_intf_1094.finish = finish;
    csv_file_dump fifo_csv_dumper_1094;
    csv_file_dump cstatus_csv_dumper_1094;
    df_fifo_monitor fifo_monitor_1094;
    df_fifo_intf fifo_intf_1095(clock,reset);
    assign fifo_intf_1095.rd_en = AESL_inst_myproject.layer2_out_1094_U.if_read & AESL_inst_myproject.layer2_out_1094_U.if_empty_n;
    assign fifo_intf_1095.wr_en = AESL_inst_myproject.layer2_out_1094_U.if_write & AESL_inst_myproject.layer2_out_1094_U.if_full_n;
    assign fifo_intf_1095.fifo_rd_block = 0;
    assign fifo_intf_1095.fifo_wr_block = 0;
    assign fifo_intf_1095.finish = finish;
    csv_file_dump fifo_csv_dumper_1095;
    csv_file_dump cstatus_csv_dumper_1095;
    df_fifo_monitor fifo_monitor_1095;
    df_fifo_intf fifo_intf_1096(clock,reset);
    assign fifo_intf_1096.rd_en = AESL_inst_myproject.layer2_out_1095_U.if_read & AESL_inst_myproject.layer2_out_1095_U.if_empty_n;
    assign fifo_intf_1096.wr_en = AESL_inst_myproject.layer2_out_1095_U.if_write & AESL_inst_myproject.layer2_out_1095_U.if_full_n;
    assign fifo_intf_1096.fifo_rd_block = 0;
    assign fifo_intf_1096.fifo_wr_block = 0;
    assign fifo_intf_1096.finish = finish;
    csv_file_dump fifo_csv_dumper_1096;
    csv_file_dump cstatus_csv_dumper_1096;
    df_fifo_monitor fifo_monitor_1096;
    df_fifo_intf fifo_intf_1097(clock,reset);
    assign fifo_intf_1097.rd_en = AESL_inst_myproject.layer2_out_1096_U.if_read & AESL_inst_myproject.layer2_out_1096_U.if_empty_n;
    assign fifo_intf_1097.wr_en = AESL_inst_myproject.layer2_out_1096_U.if_write & AESL_inst_myproject.layer2_out_1096_U.if_full_n;
    assign fifo_intf_1097.fifo_rd_block = 0;
    assign fifo_intf_1097.fifo_wr_block = 0;
    assign fifo_intf_1097.finish = finish;
    csv_file_dump fifo_csv_dumper_1097;
    csv_file_dump cstatus_csv_dumper_1097;
    df_fifo_monitor fifo_monitor_1097;
    df_fifo_intf fifo_intf_1098(clock,reset);
    assign fifo_intf_1098.rd_en = AESL_inst_myproject.layer2_out_1097_U.if_read & AESL_inst_myproject.layer2_out_1097_U.if_empty_n;
    assign fifo_intf_1098.wr_en = AESL_inst_myproject.layer2_out_1097_U.if_write & AESL_inst_myproject.layer2_out_1097_U.if_full_n;
    assign fifo_intf_1098.fifo_rd_block = 0;
    assign fifo_intf_1098.fifo_wr_block = 0;
    assign fifo_intf_1098.finish = finish;
    csv_file_dump fifo_csv_dumper_1098;
    csv_file_dump cstatus_csv_dumper_1098;
    df_fifo_monitor fifo_monitor_1098;
    df_fifo_intf fifo_intf_1099(clock,reset);
    assign fifo_intf_1099.rd_en = AESL_inst_myproject.layer2_out_1098_U.if_read & AESL_inst_myproject.layer2_out_1098_U.if_empty_n;
    assign fifo_intf_1099.wr_en = AESL_inst_myproject.layer2_out_1098_U.if_write & AESL_inst_myproject.layer2_out_1098_U.if_full_n;
    assign fifo_intf_1099.fifo_rd_block = 0;
    assign fifo_intf_1099.fifo_wr_block = 0;
    assign fifo_intf_1099.finish = finish;
    csv_file_dump fifo_csv_dumper_1099;
    csv_file_dump cstatus_csv_dumper_1099;
    df_fifo_monitor fifo_monitor_1099;
    df_fifo_intf fifo_intf_1100(clock,reset);
    assign fifo_intf_1100.rd_en = AESL_inst_myproject.layer2_out_1099_U.if_read & AESL_inst_myproject.layer2_out_1099_U.if_empty_n;
    assign fifo_intf_1100.wr_en = AESL_inst_myproject.layer2_out_1099_U.if_write & AESL_inst_myproject.layer2_out_1099_U.if_full_n;
    assign fifo_intf_1100.fifo_rd_block = 0;
    assign fifo_intf_1100.fifo_wr_block = 0;
    assign fifo_intf_1100.finish = finish;
    csv_file_dump fifo_csv_dumper_1100;
    csv_file_dump cstatus_csv_dumper_1100;
    df_fifo_monitor fifo_monitor_1100;
    df_fifo_intf fifo_intf_1101(clock,reset);
    assign fifo_intf_1101.rd_en = AESL_inst_myproject.layer2_out_1100_U.if_read & AESL_inst_myproject.layer2_out_1100_U.if_empty_n;
    assign fifo_intf_1101.wr_en = AESL_inst_myproject.layer2_out_1100_U.if_write & AESL_inst_myproject.layer2_out_1100_U.if_full_n;
    assign fifo_intf_1101.fifo_rd_block = 0;
    assign fifo_intf_1101.fifo_wr_block = 0;
    assign fifo_intf_1101.finish = finish;
    csv_file_dump fifo_csv_dumper_1101;
    csv_file_dump cstatus_csv_dumper_1101;
    df_fifo_monitor fifo_monitor_1101;
    df_fifo_intf fifo_intf_1102(clock,reset);
    assign fifo_intf_1102.rd_en = AESL_inst_myproject.layer2_out_1101_U.if_read & AESL_inst_myproject.layer2_out_1101_U.if_empty_n;
    assign fifo_intf_1102.wr_en = AESL_inst_myproject.layer2_out_1101_U.if_write & AESL_inst_myproject.layer2_out_1101_U.if_full_n;
    assign fifo_intf_1102.fifo_rd_block = 0;
    assign fifo_intf_1102.fifo_wr_block = 0;
    assign fifo_intf_1102.finish = finish;
    csv_file_dump fifo_csv_dumper_1102;
    csv_file_dump cstatus_csv_dumper_1102;
    df_fifo_monitor fifo_monitor_1102;
    df_fifo_intf fifo_intf_1103(clock,reset);
    assign fifo_intf_1103.rd_en = AESL_inst_myproject.layer2_out_1102_U.if_read & AESL_inst_myproject.layer2_out_1102_U.if_empty_n;
    assign fifo_intf_1103.wr_en = AESL_inst_myproject.layer2_out_1102_U.if_write & AESL_inst_myproject.layer2_out_1102_U.if_full_n;
    assign fifo_intf_1103.fifo_rd_block = 0;
    assign fifo_intf_1103.fifo_wr_block = 0;
    assign fifo_intf_1103.finish = finish;
    csv_file_dump fifo_csv_dumper_1103;
    csv_file_dump cstatus_csv_dumper_1103;
    df_fifo_monitor fifo_monitor_1103;
    df_fifo_intf fifo_intf_1104(clock,reset);
    assign fifo_intf_1104.rd_en = AESL_inst_myproject.layer2_out_1103_U.if_read & AESL_inst_myproject.layer2_out_1103_U.if_empty_n;
    assign fifo_intf_1104.wr_en = AESL_inst_myproject.layer2_out_1103_U.if_write & AESL_inst_myproject.layer2_out_1103_U.if_full_n;
    assign fifo_intf_1104.fifo_rd_block = 0;
    assign fifo_intf_1104.fifo_wr_block = 0;
    assign fifo_intf_1104.finish = finish;
    csv_file_dump fifo_csv_dumper_1104;
    csv_file_dump cstatus_csv_dumper_1104;
    df_fifo_monitor fifo_monitor_1104;
    df_fifo_intf fifo_intf_1105(clock,reset);
    assign fifo_intf_1105.rd_en = AESL_inst_myproject.layer2_out_1104_U.if_read & AESL_inst_myproject.layer2_out_1104_U.if_empty_n;
    assign fifo_intf_1105.wr_en = AESL_inst_myproject.layer2_out_1104_U.if_write & AESL_inst_myproject.layer2_out_1104_U.if_full_n;
    assign fifo_intf_1105.fifo_rd_block = 0;
    assign fifo_intf_1105.fifo_wr_block = 0;
    assign fifo_intf_1105.finish = finish;
    csv_file_dump fifo_csv_dumper_1105;
    csv_file_dump cstatus_csv_dumper_1105;
    df_fifo_monitor fifo_monitor_1105;
    df_fifo_intf fifo_intf_1106(clock,reset);
    assign fifo_intf_1106.rd_en = AESL_inst_myproject.layer2_out_1105_U.if_read & AESL_inst_myproject.layer2_out_1105_U.if_empty_n;
    assign fifo_intf_1106.wr_en = AESL_inst_myproject.layer2_out_1105_U.if_write & AESL_inst_myproject.layer2_out_1105_U.if_full_n;
    assign fifo_intf_1106.fifo_rd_block = 0;
    assign fifo_intf_1106.fifo_wr_block = 0;
    assign fifo_intf_1106.finish = finish;
    csv_file_dump fifo_csv_dumper_1106;
    csv_file_dump cstatus_csv_dumper_1106;
    df_fifo_monitor fifo_monitor_1106;
    df_fifo_intf fifo_intf_1107(clock,reset);
    assign fifo_intf_1107.rd_en = AESL_inst_myproject.layer2_out_1106_U.if_read & AESL_inst_myproject.layer2_out_1106_U.if_empty_n;
    assign fifo_intf_1107.wr_en = AESL_inst_myproject.layer2_out_1106_U.if_write & AESL_inst_myproject.layer2_out_1106_U.if_full_n;
    assign fifo_intf_1107.fifo_rd_block = 0;
    assign fifo_intf_1107.fifo_wr_block = 0;
    assign fifo_intf_1107.finish = finish;
    csv_file_dump fifo_csv_dumper_1107;
    csv_file_dump cstatus_csv_dumper_1107;
    df_fifo_monitor fifo_monitor_1107;
    df_fifo_intf fifo_intf_1108(clock,reset);
    assign fifo_intf_1108.rd_en = AESL_inst_myproject.layer2_out_1107_U.if_read & AESL_inst_myproject.layer2_out_1107_U.if_empty_n;
    assign fifo_intf_1108.wr_en = AESL_inst_myproject.layer2_out_1107_U.if_write & AESL_inst_myproject.layer2_out_1107_U.if_full_n;
    assign fifo_intf_1108.fifo_rd_block = 0;
    assign fifo_intf_1108.fifo_wr_block = 0;
    assign fifo_intf_1108.finish = finish;
    csv_file_dump fifo_csv_dumper_1108;
    csv_file_dump cstatus_csv_dumper_1108;
    df_fifo_monitor fifo_monitor_1108;
    df_fifo_intf fifo_intf_1109(clock,reset);
    assign fifo_intf_1109.rd_en = AESL_inst_myproject.layer2_out_1108_U.if_read & AESL_inst_myproject.layer2_out_1108_U.if_empty_n;
    assign fifo_intf_1109.wr_en = AESL_inst_myproject.layer2_out_1108_U.if_write & AESL_inst_myproject.layer2_out_1108_U.if_full_n;
    assign fifo_intf_1109.fifo_rd_block = 0;
    assign fifo_intf_1109.fifo_wr_block = 0;
    assign fifo_intf_1109.finish = finish;
    csv_file_dump fifo_csv_dumper_1109;
    csv_file_dump cstatus_csv_dumper_1109;
    df_fifo_monitor fifo_monitor_1109;
    df_fifo_intf fifo_intf_1110(clock,reset);
    assign fifo_intf_1110.rd_en = AESL_inst_myproject.layer2_out_1109_U.if_read & AESL_inst_myproject.layer2_out_1109_U.if_empty_n;
    assign fifo_intf_1110.wr_en = AESL_inst_myproject.layer2_out_1109_U.if_write & AESL_inst_myproject.layer2_out_1109_U.if_full_n;
    assign fifo_intf_1110.fifo_rd_block = 0;
    assign fifo_intf_1110.fifo_wr_block = 0;
    assign fifo_intf_1110.finish = finish;
    csv_file_dump fifo_csv_dumper_1110;
    csv_file_dump cstatus_csv_dumper_1110;
    df_fifo_monitor fifo_monitor_1110;
    df_fifo_intf fifo_intf_1111(clock,reset);
    assign fifo_intf_1111.rd_en = AESL_inst_myproject.layer2_out_1110_U.if_read & AESL_inst_myproject.layer2_out_1110_U.if_empty_n;
    assign fifo_intf_1111.wr_en = AESL_inst_myproject.layer2_out_1110_U.if_write & AESL_inst_myproject.layer2_out_1110_U.if_full_n;
    assign fifo_intf_1111.fifo_rd_block = 0;
    assign fifo_intf_1111.fifo_wr_block = 0;
    assign fifo_intf_1111.finish = finish;
    csv_file_dump fifo_csv_dumper_1111;
    csv_file_dump cstatus_csv_dumper_1111;
    df_fifo_monitor fifo_monitor_1111;
    df_fifo_intf fifo_intf_1112(clock,reset);
    assign fifo_intf_1112.rd_en = AESL_inst_myproject.layer2_out_1111_U.if_read & AESL_inst_myproject.layer2_out_1111_U.if_empty_n;
    assign fifo_intf_1112.wr_en = AESL_inst_myproject.layer2_out_1111_U.if_write & AESL_inst_myproject.layer2_out_1111_U.if_full_n;
    assign fifo_intf_1112.fifo_rd_block = 0;
    assign fifo_intf_1112.fifo_wr_block = 0;
    assign fifo_intf_1112.finish = finish;
    csv_file_dump fifo_csv_dumper_1112;
    csv_file_dump cstatus_csv_dumper_1112;
    df_fifo_monitor fifo_monitor_1112;
    df_fifo_intf fifo_intf_1113(clock,reset);
    assign fifo_intf_1113.rd_en = AESL_inst_myproject.layer2_out_1112_U.if_read & AESL_inst_myproject.layer2_out_1112_U.if_empty_n;
    assign fifo_intf_1113.wr_en = AESL_inst_myproject.layer2_out_1112_U.if_write & AESL_inst_myproject.layer2_out_1112_U.if_full_n;
    assign fifo_intf_1113.fifo_rd_block = 0;
    assign fifo_intf_1113.fifo_wr_block = 0;
    assign fifo_intf_1113.finish = finish;
    csv_file_dump fifo_csv_dumper_1113;
    csv_file_dump cstatus_csv_dumper_1113;
    df_fifo_monitor fifo_monitor_1113;
    df_fifo_intf fifo_intf_1114(clock,reset);
    assign fifo_intf_1114.rd_en = AESL_inst_myproject.layer2_out_1113_U.if_read & AESL_inst_myproject.layer2_out_1113_U.if_empty_n;
    assign fifo_intf_1114.wr_en = AESL_inst_myproject.layer2_out_1113_U.if_write & AESL_inst_myproject.layer2_out_1113_U.if_full_n;
    assign fifo_intf_1114.fifo_rd_block = 0;
    assign fifo_intf_1114.fifo_wr_block = 0;
    assign fifo_intf_1114.finish = finish;
    csv_file_dump fifo_csv_dumper_1114;
    csv_file_dump cstatus_csv_dumper_1114;
    df_fifo_monitor fifo_monitor_1114;
    df_fifo_intf fifo_intf_1115(clock,reset);
    assign fifo_intf_1115.rd_en = AESL_inst_myproject.layer2_out_1114_U.if_read & AESL_inst_myproject.layer2_out_1114_U.if_empty_n;
    assign fifo_intf_1115.wr_en = AESL_inst_myproject.layer2_out_1114_U.if_write & AESL_inst_myproject.layer2_out_1114_U.if_full_n;
    assign fifo_intf_1115.fifo_rd_block = 0;
    assign fifo_intf_1115.fifo_wr_block = 0;
    assign fifo_intf_1115.finish = finish;
    csv_file_dump fifo_csv_dumper_1115;
    csv_file_dump cstatus_csv_dumper_1115;
    df_fifo_monitor fifo_monitor_1115;
    df_fifo_intf fifo_intf_1116(clock,reset);
    assign fifo_intf_1116.rd_en = AESL_inst_myproject.layer2_out_1115_U.if_read & AESL_inst_myproject.layer2_out_1115_U.if_empty_n;
    assign fifo_intf_1116.wr_en = AESL_inst_myproject.layer2_out_1115_U.if_write & AESL_inst_myproject.layer2_out_1115_U.if_full_n;
    assign fifo_intf_1116.fifo_rd_block = 0;
    assign fifo_intf_1116.fifo_wr_block = 0;
    assign fifo_intf_1116.finish = finish;
    csv_file_dump fifo_csv_dumper_1116;
    csv_file_dump cstatus_csv_dumper_1116;
    df_fifo_monitor fifo_monitor_1116;
    df_fifo_intf fifo_intf_1117(clock,reset);
    assign fifo_intf_1117.rd_en = AESL_inst_myproject.layer2_out_1116_U.if_read & AESL_inst_myproject.layer2_out_1116_U.if_empty_n;
    assign fifo_intf_1117.wr_en = AESL_inst_myproject.layer2_out_1116_U.if_write & AESL_inst_myproject.layer2_out_1116_U.if_full_n;
    assign fifo_intf_1117.fifo_rd_block = 0;
    assign fifo_intf_1117.fifo_wr_block = 0;
    assign fifo_intf_1117.finish = finish;
    csv_file_dump fifo_csv_dumper_1117;
    csv_file_dump cstatus_csv_dumper_1117;
    df_fifo_monitor fifo_monitor_1117;
    df_fifo_intf fifo_intf_1118(clock,reset);
    assign fifo_intf_1118.rd_en = AESL_inst_myproject.layer2_out_1117_U.if_read & AESL_inst_myproject.layer2_out_1117_U.if_empty_n;
    assign fifo_intf_1118.wr_en = AESL_inst_myproject.layer2_out_1117_U.if_write & AESL_inst_myproject.layer2_out_1117_U.if_full_n;
    assign fifo_intf_1118.fifo_rd_block = 0;
    assign fifo_intf_1118.fifo_wr_block = 0;
    assign fifo_intf_1118.finish = finish;
    csv_file_dump fifo_csv_dumper_1118;
    csv_file_dump cstatus_csv_dumper_1118;
    df_fifo_monitor fifo_monitor_1118;
    df_fifo_intf fifo_intf_1119(clock,reset);
    assign fifo_intf_1119.rd_en = AESL_inst_myproject.layer2_out_1118_U.if_read & AESL_inst_myproject.layer2_out_1118_U.if_empty_n;
    assign fifo_intf_1119.wr_en = AESL_inst_myproject.layer2_out_1118_U.if_write & AESL_inst_myproject.layer2_out_1118_U.if_full_n;
    assign fifo_intf_1119.fifo_rd_block = 0;
    assign fifo_intf_1119.fifo_wr_block = 0;
    assign fifo_intf_1119.finish = finish;
    csv_file_dump fifo_csv_dumper_1119;
    csv_file_dump cstatus_csv_dumper_1119;
    df_fifo_monitor fifo_monitor_1119;
    df_fifo_intf fifo_intf_1120(clock,reset);
    assign fifo_intf_1120.rd_en = AESL_inst_myproject.layer2_out_1119_U.if_read & AESL_inst_myproject.layer2_out_1119_U.if_empty_n;
    assign fifo_intf_1120.wr_en = AESL_inst_myproject.layer2_out_1119_U.if_write & AESL_inst_myproject.layer2_out_1119_U.if_full_n;
    assign fifo_intf_1120.fifo_rd_block = 0;
    assign fifo_intf_1120.fifo_wr_block = 0;
    assign fifo_intf_1120.finish = finish;
    csv_file_dump fifo_csv_dumper_1120;
    csv_file_dump cstatus_csv_dumper_1120;
    df_fifo_monitor fifo_monitor_1120;
    df_fifo_intf fifo_intf_1121(clock,reset);
    assign fifo_intf_1121.rd_en = AESL_inst_myproject.layer2_out_1120_U.if_read & AESL_inst_myproject.layer2_out_1120_U.if_empty_n;
    assign fifo_intf_1121.wr_en = AESL_inst_myproject.layer2_out_1120_U.if_write & AESL_inst_myproject.layer2_out_1120_U.if_full_n;
    assign fifo_intf_1121.fifo_rd_block = 0;
    assign fifo_intf_1121.fifo_wr_block = 0;
    assign fifo_intf_1121.finish = finish;
    csv_file_dump fifo_csv_dumper_1121;
    csv_file_dump cstatus_csv_dumper_1121;
    df_fifo_monitor fifo_monitor_1121;
    df_fifo_intf fifo_intf_1122(clock,reset);
    assign fifo_intf_1122.rd_en = AESL_inst_myproject.layer2_out_1121_U.if_read & AESL_inst_myproject.layer2_out_1121_U.if_empty_n;
    assign fifo_intf_1122.wr_en = AESL_inst_myproject.layer2_out_1121_U.if_write & AESL_inst_myproject.layer2_out_1121_U.if_full_n;
    assign fifo_intf_1122.fifo_rd_block = 0;
    assign fifo_intf_1122.fifo_wr_block = 0;
    assign fifo_intf_1122.finish = finish;
    csv_file_dump fifo_csv_dumper_1122;
    csv_file_dump cstatus_csv_dumper_1122;
    df_fifo_monitor fifo_monitor_1122;
    df_fifo_intf fifo_intf_1123(clock,reset);
    assign fifo_intf_1123.rd_en = AESL_inst_myproject.layer2_out_1122_U.if_read & AESL_inst_myproject.layer2_out_1122_U.if_empty_n;
    assign fifo_intf_1123.wr_en = AESL_inst_myproject.layer2_out_1122_U.if_write & AESL_inst_myproject.layer2_out_1122_U.if_full_n;
    assign fifo_intf_1123.fifo_rd_block = 0;
    assign fifo_intf_1123.fifo_wr_block = 0;
    assign fifo_intf_1123.finish = finish;
    csv_file_dump fifo_csv_dumper_1123;
    csv_file_dump cstatus_csv_dumper_1123;
    df_fifo_monitor fifo_monitor_1123;
    df_fifo_intf fifo_intf_1124(clock,reset);
    assign fifo_intf_1124.rd_en = AESL_inst_myproject.layer2_out_1123_U.if_read & AESL_inst_myproject.layer2_out_1123_U.if_empty_n;
    assign fifo_intf_1124.wr_en = AESL_inst_myproject.layer2_out_1123_U.if_write & AESL_inst_myproject.layer2_out_1123_U.if_full_n;
    assign fifo_intf_1124.fifo_rd_block = 0;
    assign fifo_intf_1124.fifo_wr_block = 0;
    assign fifo_intf_1124.finish = finish;
    csv_file_dump fifo_csv_dumper_1124;
    csv_file_dump cstatus_csv_dumper_1124;
    df_fifo_monitor fifo_monitor_1124;
    df_fifo_intf fifo_intf_1125(clock,reset);
    assign fifo_intf_1125.rd_en = AESL_inst_myproject.layer2_out_1124_U.if_read & AESL_inst_myproject.layer2_out_1124_U.if_empty_n;
    assign fifo_intf_1125.wr_en = AESL_inst_myproject.layer2_out_1124_U.if_write & AESL_inst_myproject.layer2_out_1124_U.if_full_n;
    assign fifo_intf_1125.fifo_rd_block = 0;
    assign fifo_intf_1125.fifo_wr_block = 0;
    assign fifo_intf_1125.finish = finish;
    csv_file_dump fifo_csv_dumper_1125;
    csv_file_dump cstatus_csv_dumper_1125;
    df_fifo_monitor fifo_monitor_1125;
    df_fifo_intf fifo_intf_1126(clock,reset);
    assign fifo_intf_1126.rd_en = AESL_inst_myproject.layer2_out_1125_U.if_read & AESL_inst_myproject.layer2_out_1125_U.if_empty_n;
    assign fifo_intf_1126.wr_en = AESL_inst_myproject.layer2_out_1125_U.if_write & AESL_inst_myproject.layer2_out_1125_U.if_full_n;
    assign fifo_intf_1126.fifo_rd_block = 0;
    assign fifo_intf_1126.fifo_wr_block = 0;
    assign fifo_intf_1126.finish = finish;
    csv_file_dump fifo_csv_dumper_1126;
    csv_file_dump cstatus_csv_dumper_1126;
    df_fifo_monitor fifo_monitor_1126;
    df_fifo_intf fifo_intf_1127(clock,reset);
    assign fifo_intf_1127.rd_en = AESL_inst_myproject.layer2_out_1126_U.if_read & AESL_inst_myproject.layer2_out_1126_U.if_empty_n;
    assign fifo_intf_1127.wr_en = AESL_inst_myproject.layer2_out_1126_U.if_write & AESL_inst_myproject.layer2_out_1126_U.if_full_n;
    assign fifo_intf_1127.fifo_rd_block = 0;
    assign fifo_intf_1127.fifo_wr_block = 0;
    assign fifo_intf_1127.finish = finish;
    csv_file_dump fifo_csv_dumper_1127;
    csv_file_dump cstatus_csv_dumper_1127;
    df_fifo_monitor fifo_monitor_1127;
    df_fifo_intf fifo_intf_1128(clock,reset);
    assign fifo_intf_1128.rd_en = AESL_inst_myproject.layer2_out_1127_U.if_read & AESL_inst_myproject.layer2_out_1127_U.if_empty_n;
    assign fifo_intf_1128.wr_en = AESL_inst_myproject.layer2_out_1127_U.if_write & AESL_inst_myproject.layer2_out_1127_U.if_full_n;
    assign fifo_intf_1128.fifo_rd_block = 0;
    assign fifo_intf_1128.fifo_wr_block = 0;
    assign fifo_intf_1128.finish = finish;
    csv_file_dump fifo_csv_dumper_1128;
    csv_file_dump cstatus_csv_dumper_1128;
    df_fifo_monitor fifo_monitor_1128;
    df_fifo_intf fifo_intf_1129(clock,reset);
    assign fifo_intf_1129.rd_en = AESL_inst_myproject.layer2_out_1128_U.if_read & AESL_inst_myproject.layer2_out_1128_U.if_empty_n;
    assign fifo_intf_1129.wr_en = AESL_inst_myproject.layer2_out_1128_U.if_write & AESL_inst_myproject.layer2_out_1128_U.if_full_n;
    assign fifo_intf_1129.fifo_rd_block = 0;
    assign fifo_intf_1129.fifo_wr_block = 0;
    assign fifo_intf_1129.finish = finish;
    csv_file_dump fifo_csv_dumper_1129;
    csv_file_dump cstatus_csv_dumper_1129;
    df_fifo_monitor fifo_monitor_1129;
    df_fifo_intf fifo_intf_1130(clock,reset);
    assign fifo_intf_1130.rd_en = AESL_inst_myproject.layer2_out_1129_U.if_read & AESL_inst_myproject.layer2_out_1129_U.if_empty_n;
    assign fifo_intf_1130.wr_en = AESL_inst_myproject.layer2_out_1129_U.if_write & AESL_inst_myproject.layer2_out_1129_U.if_full_n;
    assign fifo_intf_1130.fifo_rd_block = 0;
    assign fifo_intf_1130.fifo_wr_block = 0;
    assign fifo_intf_1130.finish = finish;
    csv_file_dump fifo_csv_dumper_1130;
    csv_file_dump cstatus_csv_dumper_1130;
    df_fifo_monitor fifo_monitor_1130;
    df_fifo_intf fifo_intf_1131(clock,reset);
    assign fifo_intf_1131.rd_en = AESL_inst_myproject.layer2_out_1130_U.if_read & AESL_inst_myproject.layer2_out_1130_U.if_empty_n;
    assign fifo_intf_1131.wr_en = AESL_inst_myproject.layer2_out_1130_U.if_write & AESL_inst_myproject.layer2_out_1130_U.if_full_n;
    assign fifo_intf_1131.fifo_rd_block = 0;
    assign fifo_intf_1131.fifo_wr_block = 0;
    assign fifo_intf_1131.finish = finish;
    csv_file_dump fifo_csv_dumper_1131;
    csv_file_dump cstatus_csv_dumper_1131;
    df_fifo_monitor fifo_monitor_1131;
    df_fifo_intf fifo_intf_1132(clock,reset);
    assign fifo_intf_1132.rd_en = AESL_inst_myproject.layer2_out_1131_U.if_read & AESL_inst_myproject.layer2_out_1131_U.if_empty_n;
    assign fifo_intf_1132.wr_en = AESL_inst_myproject.layer2_out_1131_U.if_write & AESL_inst_myproject.layer2_out_1131_U.if_full_n;
    assign fifo_intf_1132.fifo_rd_block = 0;
    assign fifo_intf_1132.fifo_wr_block = 0;
    assign fifo_intf_1132.finish = finish;
    csv_file_dump fifo_csv_dumper_1132;
    csv_file_dump cstatus_csv_dumper_1132;
    df_fifo_monitor fifo_monitor_1132;
    df_fifo_intf fifo_intf_1133(clock,reset);
    assign fifo_intf_1133.rd_en = AESL_inst_myproject.layer2_out_1132_U.if_read & AESL_inst_myproject.layer2_out_1132_U.if_empty_n;
    assign fifo_intf_1133.wr_en = AESL_inst_myproject.layer2_out_1132_U.if_write & AESL_inst_myproject.layer2_out_1132_U.if_full_n;
    assign fifo_intf_1133.fifo_rd_block = 0;
    assign fifo_intf_1133.fifo_wr_block = 0;
    assign fifo_intf_1133.finish = finish;
    csv_file_dump fifo_csv_dumper_1133;
    csv_file_dump cstatus_csv_dumper_1133;
    df_fifo_monitor fifo_monitor_1133;
    df_fifo_intf fifo_intf_1134(clock,reset);
    assign fifo_intf_1134.rd_en = AESL_inst_myproject.layer2_out_1133_U.if_read & AESL_inst_myproject.layer2_out_1133_U.if_empty_n;
    assign fifo_intf_1134.wr_en = AESL_inst_myproject.layer2_out_1133_U.if_write & AESL_inst_myproject.layer2_out_1133_U.if_full_n;
    assign fifo_intf_1134.fifo_rd_block = 0;
    assign fifo_intf_1134.fifo_wr_block = 0;
    assign fifo_intf_1134.finish = finish;
    csv_file_dump fifo_csv_dumper_1134;
    csv_file_dump cstatus_csv_dumper_1134;
    df_fifo_monitor fifo_monitor_1134;
    df_fifo_intf fifo_intf_1135(clock,reset);
    assign fifo_intf_1135.rd_en = AESL_inst_myproject.layer2_out_1134_U.if_read & AESL_inst_myproject.layer2_out_1134_U.if_empty_n;
    assign fifo_intf_1135.wr_en = AESL_inst_myproject.layer2_out_1134_U.if_write & AESL_inst_myproject.layer2_out_1134_U.if_full_n;
    assign fifo_intf_1135.fifo_rd_block = 0;
    assign fifo_intf_1135.fifo_wr_block = 0;
    assign fifo_intf_1135.finish = finish;
    csv_file_dump fifo_csv_dumper_1135;
    csv_file_dump cstatus_csv_dumper_1135;
    df_fifo_monitor fifo_monitor_1135;
    df_fifo_intf fifo_intf_1136(clock,reset);
    assign fifo_intf_1136.rd_en = AESL_inst_myproject.layer2_out_1135_U.if_read & AESL_inst_myproject.layer2_out_1135_U.if_empty_n;
    assign fifo_intf_1136.wr_en = AESL_inst_myproject.layer2_out_1135_U.if_write & AESL_inst_myproject.layer2_out_1135_U.if_full_n;
    assign fifo_intf_1136.fifo_rd_block = 0;
    assign fifo_intf_1136.fifo_wr_block = 0;
    assign fifo_intf_1136.finish = finish;
    csv_file_dump fifo_csv_dumper_1136;
    csv_file_dump cstatus_csv_dumper_1136;
    df_fifo_monitor fifo_monitor_1136;
    df_fifo_intf fifo_intf_1137(clock,reset);
    assign fifo_intf_1137.rd_en = AESL_inst_myproject.layer2_out_1136_U.if_read & AESL_inst_myproject.layer2_out_1136_U.if_empty_n;
    assign fifo_intf_1137.wr_en = AESL_inst_myproject.layer2_out_1136_U.if_write & AESL_inst_myproject.layer2_out_1136_U.if_full_n;
    assign fifo_intf_1137.fifo_rd_block = 0;
    assign fifo_intf_1137.fifo_wr_block = 0;
    assign fifo_intf_1137.finish = finish;
    csv_file_dump fifo_csv_dumper_1137;
    csv_file_dump cstatus_csv_dumper_1137;
    df_fifo_monitor fifo_monitor_1137;
    df_fifo_intf fifo_intf_1138(clock,reset);
    assign fifo_intf_1138.rd_en = AESL_inst_myproject.layer2_out_1137_U.if_read & AESL_inst_myproject.layer2_out_1137_U.if_empty_n;
    assign fifo_intf_1138.wr_en = AESL_inst_myproject.layer2_out_1137_U.if_write & AESL_inst_myproject.layer2_out_1137_U.if_full_n;
    assign fifo_intf_1138.fifo_rd_block = 0;
    assign fifo_intf_1138.fifo_wr_block = 0;
    assign fifo_intf_1138.finish = finish;
    csv_file_dump fifo_csv_dumper_1138;
    csv_file_dump cstatus_csv_dumper_1138;
    df_fifo_monitor fifo_monitor_1138;
    df_fifo_intf fifo_intf_1139(clock,reset);
    assign fifo_intf_1139.rd_en = AESL_inst_myproject.layer2_out_1138_U.if_read & AESL_inst_myproject.layer2_out_1138_U.if_empty_n;
    assign fifo_intf_1139.wr_en = AESL_inst_myproject.layer2_out_1138_U.if_write & AESL_inst_myproject.layer2_out_1138_U.if_full_n;
    assign fifo_intf_1139.fifo_rd_block = 0;
    assign fifo_intf_1139.fifo_wr_block = 0;
    assign fifo_intf_1139.finish = finish;
    csv_file_dump fifo_csv_dumper_1139;
    csv_file_dump cstatus_csv_dumper_1139;
    df_fifo_monitor fifo_monitor_1139;
    df_fifo_intf fifo_intf_1140(clock,reset);
    assign fifo_intf_1140.rd_en = AESL_inst_myproject.layer2_out_1139_U.if_read & AESL_inst_myproject.layer2_out_1139_U.if_empty_n;
    assign fifo_intf_1140.wr_en = AESL_inst_myproject.layer2_out_1139_U.if_write & AESL_inst_myproject.layer2_out_1139_U.if_full_n;
    assign fifo_intf_1140.fifo_rd_block = 0;
    assign fifo_intf_1140.fifo_wr_block = 0;
    assign fifo_intf_1140.finish = finish;
    csv_file_dump fifo_csv_dumper_1140;
    csv_file_dump cstatus_csv_dumper_1140;
    df_fifo_monitor fifo_monitor_1140;
    df_fifo_intf fifo_intf_1141(clock,reset);
    assign fifo_intf_1141.rd_en = AESL_inst_myproject.layer2_out_1140_U.if_read & AESL_inst_myproject.layer2_out_1140_U.if_empty_n;
    assign fifo_intf_1141.wr_en = AESL_inst_myproject.layer2_out_1140_U.if_write & AESL_inst_myproject.layer2_out_1140_U.if_full_n;
    assign fifo_intf_1141.fifo_rd_block = 0;
    assign fifo_intf_1141.fifo_wr_block = 0;
    assign fifo_intf_1141.finish = finish;
    csv_file_dump fifo_csv_dumper_1141;
    csv_file_dump cstatus_csv_dumper_1141;
    df_fifo_monitor fifo_monitor_1141;
    df_fifo_intf fifo_intf_1142(clock,reset);
    assign fifo_intf_1142.rd_en = AESL_inst_myproject.layer2_out_1141_U.if_read & AESL_inst_myproject.layer2_out_1141_U.if_empty_n;
    assign fifo_intf_1142.wr_en = AESL_inst_myproject.layer2_out_1141_U.if_write & AESL_inst_myproject.layer2_out_1141_U.if_full_n;
    assign fifo_intf_1142.fifo_rd_block = 0;
    assign fifo_intf_1142.fifo_wr_block = 0;
    assign fifo_intf_1142.finish = finish;
    csv_file_dump fifo_csv_dumper_1142;
    csv_file_dump cstatus_csv_dumper_1142;
    df_fifo_monitor fifo_monitor_1142;
    df_fifo_intf fifo_intf_1143(clock,reset);
    assign fifo_intf_1143.rd_en = AESL_inst_myproject.layer2_out_1142_U.if_read & AESL_inst_myproject.layer2_out_1142_U.if_empty_n;
    assign fifo_intf_1143.wr_en = AESL_inst_myproject.layer2_out_1142_U.if_write & AESL_inst_myproject.layer2_out_1142_U.if_full_n;
    assign fifo_intf_1143.fifo_rd_block = 0;
    assign fifo_intf_1143.fifo_wr_block = 0;
    assign fifo_intf_1143.finish = finish;
    csv_file_dump fifo_csv_dumper_1143;
    csv_file_dump cstatus_csv_dumper_1143;
    df_fifo_monitor fifo_monitor_1143;
    df_fifo_intf fifo_intf_1144(clock,reset);
    assign fifo_intf_1144.rd_en = AESL_inst_myproject.layer2_out_1143_U.if_read & AESL_inst_myproject.layer2_out_1143_U.if_empty_n;
    assign fifo_intf_1144.wr_en = AESL_inst_myproject.layer2_out_1143_U.if_write & AESL_inst_myproject.layer2_out_1143_U.if_full_n;
    assign fifo_intf_1144.fifo_rd_block = 0;
    assign fifo_intf_1144.fifo_wr_block = 0;
    assign fifo_intf_1144.finish = finish;
    csv_file_dump fifo_csv_dumper_1144;
    csv_file_dump cstatus_csv_dumper_1144;
    df_fifo_monitor fifo_monitor_1144;
    df_fifo_intf fifo_intf_1145(clock,reset);
    assign fifo_intf_1145.rd_en = AESL_inst_myproject.layer2_out_1144_U.if_read & AESL_inst_myproject.layer2_out_1144_U.if_empty_n;
    assign fifo_intf_1145.wr_en = AESL_inst_myproject.layer2_out_1144_U.if_write & AESL_inst_myproject.layer2_out_1144_U.if_full_n;
    assign fifo_intf_1145.fifo_rd_block = 0;
    assign fifo_intf_1145.fifo_wr_block = 0;
    assign fifo_intf_1145.finish = finish;
    csv_file_dump fifo_csv_dumper_1145;
    csv_file_dump cstatus_csv_dumper_1145;
    df_fifo_monitor fifo_monitor_1145;
    df_fifo_intf fifo_intf_1146(clock,reset);
    assign fifo_intf_1146.rd_en = AESL_inst_myproject.layer2_out_1145_U.if_read & AESL_inst_myproject.layer2_out_1145_U.if_empty_n;
    assign fifo_intf_1146.wr_en = AESL_inst_myproject.layer2_out_1145_U.if_write & AESL_inst_myproject.layer2_out_1145_U.if_full_n;
    assign fifo_intf_1146.fifo_rd_block = 0;
    assign fifo_intf_1146.fifo_wr_block = 0;
    assign fifo_intf_1146.finish = finish;
    csv_file_dump fifo_csv_dumper_1146;
    csv_file_dump cstatus_csv_dumper_1146;
    df_fifo_monitor fifo_monitor_1146;
    df_fifo_intf fifo_intf_1147(clock,reset);
    assign fifo_intf_1147.rd_en = AESL_inst_myproject.layer2_out_1146_U.if_read & AESL_inst_myproject.layer2_out_1146_U.if_empty_n;
    assign fifo_intf_1147.wr_en = AESL_inst_myproject.layer2_out_1146_U.if_write & AESL_inst_myproject.layer2_out_1146_U.if_full_n;
    assign fifo_intf_1147.fifo_rd_block = 0;
    assign fifo_intf_1147.fifo_wr_block = 0;
    assign fifo_intf_1147.finish = finish;
    csv_file_dump fifo_csv_dumper_1147;
    csv_file_dump cstatus_csv_dumper_1147;
    df_fifo_monitor fifo_monitor_1147;
    df_fifo_intf fifo_intf_1148(clock,reset);
    assign fifo_intf_1148.rd_en = AESL_inst_myproject.layer2_out_1147_U.if_read & AESL_inst_myproject.layer2_out_1147_U.if_empty_n;
    assign fifo_intf_1148.wr_en = AESL_inst_myproject.layer2_out_1147_U.if_write & AESL_inst_myproject.layer2_out_1147_U.if_full_n;
    assign fifo_intf_1148.fifo_rd_block = 0;
    assign fifo_intf_1148.fifo_wr_block = 0;
    assign fifo_intf_1148.finish = finish;
    csv_file_dump fifo_csv_dumper_1148;
    csv_file_dump cstatus_csv_dumper_1148;
    df_fifo_monitor fifo_monitor_1148;
    df_fifo_intf fifo_intf_1149(clock,reset);
    assign fifo_intf_1149.rd_en = AESL_inst_myproject.layer2_out_1148_U.if_read & AESL_inst_myproject.layer2_out_1148_U.if_empty_n;
    assign fifo_intf_1149.wr_en = AESL_inst_myproject.layer2_out_1148_U.if_write & AESL_inst_myproject.layer2_out_1148_U.if_full_n;
    assign fifo_intf_1149.fifo_rd_block = 0;
    assign fifo_intf_1149.fifo_wr_block = 0;
    assign fifo_intf_1149.finish = finish;
    csv_file_dump fifo_csv_dumper_1149;
    csv_file_dump cstatus_csv_dumper_1149;
    df_fifo_monitor fifo_monitor_1149;
    df_fifo_intf fifo_intf_1150(clock,reset);
    assign fifo_intf_1150.rd_en = AESL_inst_myproject.layer2_out_1149_U.if_read & AESL_inst_myproject.layer2_out_1149_U.if_empty_n;
    assign fifo_intf_1150.wr_en = AESL_inst_myproject.layer2_out_1149_U.if_write & AESL_inst_myproject.layer2_out_1149_U.if_full_n;
    assign fifo_intf_1150.fifo_rd_block = 0;
    assign fifo_intf_1150.fifo_wr_block = 0;
    assign fifo_intf_1150.finish = finish;
    csv_file_dump fifo_csv_dumper_1150;
    csv_file_dump cstatus_csv_dumper_1150;
    df_fifo_monitor fifo_monitor_1150;
    df_fifo_intf fifo_intf_1151(clock,reset);
    assign fifo_intf_1151.rd_en = AESL_inst_myproject.layer2_out_1150_U.if_read & AESL_inst_myproject.layer2_out_1150_U.if_empty_n;
    assign fifo_intf_1151.wr_en = AESL_inst_myproject.layer2_out_1150_U.if_write & AESL_inst_myproject.layer2_out_1150_U.if_full_n;
    assign fifo_intf_1151.fifo_rd_block = 0;
    assign fifo_intf_1151.fifo_wr_block = 0;
    assign fifo_intf_1151.finish = finish;
    csv_file_dump fifo_csv_dumper_1151;
    csv_file_dump cstatus_csv_dumper_1151;
    df_fifo_monitor fifo_monitor_1151;
    df_fifo_intf fifo_intf_1152(clock,reset);
    assign fifo_intf_1152.rd_en = AESL_inst_myproject.layer2_out_1151_U.if_read & AESL_inst_myproject.layer2_out_1151_U.if_empty_n;
    assign fifo_intf_1152.wr_en = AESL_inst_myproject.layer2_out_1151_U.if_write & AESL_inst_myproject.layer2_out_1151_U.if_full_n;
    assign fifo_intf_1152.fifo_rd_block = 0;
    assign fifo_intf_1152.fifo_wr_block = 0;
    assign fifo_intf_1152.finish = finish;
    csv_file_dump fifo_csv_dumper_1152;
    csv_file_dump cstatus_csv_dumper_1152;
    df_fifo_monitor fifo_monitor_1152;
    df_fifo_intf fifo_intf_1153(clock,reset);
    assign fifo_intf_1153.rd_en = AESL_inst_myproject.layer2_out_1152_U.if_read & AESL_inst_myproject.layer2_out_1152_U.if_empty_n;
    assign fifo_intf_1153.wr_en = AESL_inst_myproject.layer2_out_1152_U.if_write & AESL_inst_myproject.layer2_out_1152_U.if_full_n;
    assign fifo_intf_1153.fifo_rd_block = 0;
    assign fifo_intf_1153.fifo_wr_block = 0;
    assign fifo_intf_1153.finish = finish;
    csv_file_dump fifo_csv_dumper_1153;
    csv_file_dump cstatus_csv_dumper_1153;
    df_fifo_monitor fifo_monitor_1153;
    df_fifo_intf fifo_intf_1154(clock,reset);
    assign fifo_intf_1154.rd_en = AESL_inst_myproject.layer2_out_1153_U.if_read & AESL_inst_myproject.layer2_out_1153_U.if_empty_n;
    assign fifo_intf_1154.wr_en = AESL_inst_myproject.layer2_out_1153_U.if_write & AESL_inst_myproject.layer2_out_1153_U.if_full_n;
    assign fifo_intf_1154.fifo_rd_block = 0;
    assign fifo_intf_1154.fifo_wr_block = 0;
    assign fifo_intf_1154.finish = finish;
    csv_file_dump fifo_csv_dumper_1154;
    csv_file_dump cstatus_csv_dumper_1154;
    df_fifo_monitor fifo_monitor_1154;
    df_fifo_intf fifo_intf_1155(clock,reset);
    assign fifo_intf_1155.rd_en = AESL_inst_myproject.layer2_out_1154_U.if_read & AESL_inst_myproject.layer2_out_1154_U.if_empty_n;
    assign fifo_intf_1155.wr_en = AESL_inst_myproject.layer2_out_1154_U.if_write & AESL_inst_myproject.layer2_out_1154_U.if_full_n;
    assign fifo_intf_1155.fifo_rd_block = 0;
    assign fifo_intf_1155.fifo_wr_block = 0;
    assign fifo_intf_1155.finish = finish;
    csv_file_dump fifo_csv_dumper_1155;
    csv_file_dump cstatus_csv_dumper_1155;
    df_fifo_monitor fifo_monitor_1155;
    df_fifo_intf fifo_intf_1156(clock,reset);
    assign fifo_intf_1156.rd_en = AESL_inst_myproject.layer2_out_1155_U.if_read & AESL_inst_myproject.layer2_out_1155_U.if_empty_n;
    assign fifo_intf_1156.wr_en = AESL_inst_myproject.layer2_out_1155_U.if_write & AESL_inst_myproject.layer2_out_1155_U.if_full_n;
    assign fifo_intf_1156.fifo_rd_block = 0;
    assign fifo_intf_1156.fifo_wr_block = 0;
    assign fifo_intf_1156.finish = finish;
    csv_file_dump fifo_csv_dumper_1156;
    csv_file_dump cstatus_csv_dumper_1156;
    df_fifo_monitor fifo_monitor_1156;
    df_fifo_intf fifo_intf_1157(clock,reset);
    assign fifo_intf_1157.rd_en = AESL_inst_myproject.layer2_out_1156_U.if_read & AESL_inst_myproject.layer2_out_1156_U.if_empty_n;
    assign fifo_intf_1157.wr_en = AESL_inst_myproject.layer2_out_1156_U.if_write & AESL_inst_myproject.layer2_out_1156_U.if_full_n;
    assign fifo_intf_1157.fifo_rd_block = 0;
    assign fifo_intf_1157.fifo_wr_block = 0;
    assign fifo_intf_1157.finish = finish;
    csv_file_dump fifo_csv_dumper_1157;
    csv_file_dump cstatus_csv_dumper_1157;
    df_fifo_monitor fifo_monitor_1157;
    df_fifo_intf fifo_intf_1158(clock,reset);
    assign fifo_intf_1158.rd_en = AESL_inst_myproject.layer2_out_1157_U.if_read & AESL_inst_myproject.layer2_out_1157_U.if_empty_n;
    assign fifo_intf_1158.wr_en = AESL_inst_myproject.layer2_out_1157_U.if_write & AESL_inst_myproject.layer2_out_1157_U.if_full_n;
    assign fifo_intf_1158.fifo_rd_block = 0;
    assign fifo_intf_1158.fifo_wr_block = 0;
    assign fifo_intf_1158.finish = finish;
    csv_file_dump fifo_csv_dumper_1158;
    csv_file_dump cstatus_csv_dumper_1158;
    df_fifo_monitor fifo_monitor_1158;
    df_fifo_intf fifo_intf_1159(clock,reset);
    assign fifo_intf_1159.rd_en = AESL_inst_myproject.layer2_out_1158_U.if_read & AESL_inst_myproject.layer2_out_1158_U.if_empty_n;
    assign fifo_intf_1159.wr_en = AESL_inst_myproject.layer2_out_1158_U.if_write & AESL_inst_myproject.layer2_out_1158_U.if_full_n;
    assign fifo_intf_1159.fifo_rd_block = 0;
    assign fifo_intf_1159.fifo_wr_block = 0;
    assign fifo_intf_1159.finish = finish;
    csv_file_dump fifo_csv_dumper_1159;
    csv_file_dump cstatus_csv_dumper_1159;
    df_fifo_monitor fifo_monitor_1159;
    df_fifo_intf fifo_intf_1160(clock,reset);
    assign fifo_intf_1160.rd_en = AESL_inst_myproject.layer2_out_1159_U.if_read & AESL_inst_myproject.layer2_out_1159_U.if_empty_n;
    assign fifo_intf_1160.wr_en = AESL_inst_myproject.layer2_out_1159_U.if_write & AESL_inst_myproject.layer2_out_1159_U.if_full_n;
    assign fifo_intf_1160.fifo_rd_block = 0;
    assign fifo_intf_1160.fifo_wr_block = 0;
    assign fifo_intf_1160.finish = finish;
    csv_file_dump fifo_csv_dumper_1160;
    csv_file_dump cstatus_csv_dumper_1160;
    df_fifo_monitor fifo_monitor_1160;
    df_fifo_intf fifo_intf_1161(clock,reset);
    assign fifo_intf_1161.rd_en = AESL_inst_myproject.layer2_out_1160_U.if_read & AESL_inst_myproject.layer2_out_1160_U.if_empty_n;
    assign fifo_intf_1161.wr_en = AESL_inst_myproject.layer2_out_1160_U.if_write & AESL_inst_myproject.layer2_out_1160_U.if_full_n;
    assign fifo_intf_1161.fifo_rd_block = 0;
    assign fifo_intf_1161.fifo_wr_block = 0;
    assign fifo_intf_1161.finish = finish;
    csv_file_dump fifo_csv_dumper_1161;
    csv_file_dump cstatus_csv_dumper_1161;
    df_fifo_monitor fifo_monitor_1161;
    df_fifo_intf fifo_intf_1162(clock,reset);
    assign fifo_intf_1162.rd_en = AESL_inst_myproject.layer2_out_1161_U.if_read & AESL_inst_myproject.layer2_out_1161_U.if_empty_n;
    assign fifo_intf_1162.wr_en = AESL_inst_myproject.layer2_out_1161_U.if_write & AESL_inst_myproject.layer2_out_1161_U.if_full_n;
    assign fifo_intf_1162.fifo_rd_block = 0;
    assign fifo_intf_1162.fifo_wr_block = 0;
    assign fifo_intf_1162.finish = finish;
    csv_file_dump fifo_csv_dumper_1162;
    csv_file_dump cstatus_csv_dumper_1162;
    df_fifo_monitor fifo_monitor_1162;
    df_fifo_intf fifo_intf_1163(clock,reset);
    assign fifo_intf_1163.rd_en = AESL_inst_myproject.layer2_out_1162_U.if_read & AESL_inst_myproject.layer2_out_1162_U.if_empty_n;
    assign fifo_intf_1163.wr_en = AESL_inst_myproject.layer2_out_1162_U.if_write & AESL_inst_myproject.layer2_out_1162_U.if_full_n;
    assign fifo_intf_1163.fifo_rd_block = 0;
    assign fifo_intf_1163.fifo_wr_block = 0;
    assign fifo_intf_1163.finish = finish;
    csv_file_dump fifo_csv_dumper_1163;
    csv_file_dump cstatus_csv_dumper_1163;
    df_fifo_monitor fifo_monitor_1163;
    df_fifo_intf fifo_intf_1164(clock,reset);
    assign fifo_intf_1164.rd_en = AESL_inst_myproject.layer2_out_1163_U.if_read & AESL_inst_myproject.layer2_out_1163_U.if_empty_n;
    assign fifo_intf_1164.wr_en = AESL_inst_myproject.layer2_out_1163_U.if_write & AESL_inst_myproject.layer2_out_1163_U.if_full_n;
    assign fifo_intf_1164.fifo_rd_block = 0;
    assign fifo_intf_1164.fifo_wr_block = 0;
    assign fifo_intf_1164.finish = finish;
    csv_file_dump fifo_csv_dumper_1164;
    csv_file_dump cstatus_csv_dumper_1164;
    df_fifo_monitor fifo_monitor_1164;
    df_fifo_intf fifo_intf_1165(clock,reset);
    assign fifo_intf_1165.rd_en = AESL_inst_myproject.layer2_out_1164_U.if_read & AESL_inst_myproject.layer2_out_1164_U.if_empty_n;
    assign fifo_intf_1165.wr_en = AESL_inst_myproject.layer2_out_1164_U.if_write & AESL_inst_myproject.layer2_out_1164_U.if_full_n;
    assign fifo_intf_1165.fifo_rd_block = 0;
    assign fifo_intf_1165.fifo_wr_block = 0;
    assign fifo_intf_1165.finish = finish;
    csv_file_dump fifo_csv_dumper_1165;
    csv_file_dump cstatus_csv_dumper_1165;
    df_fifo_monitor fifo_monitor_1165;
    df_fifo_intf fifo_intf_1166(clock,reset);
    assign fifo_intf_1166.rd_en = AESL_inst_myproject.layer2_out_1165_U.if_read & AESL_inst_myproject.layer2_out_1165_U.if_empty_n;
    assign fifo_intf_1166.wr_en = AESL_inst_myproject.layer2_out_1165_U.if_write & AESL_inst_myproject.layer2_out_1165_U.if_full_n;
    assign fifo_intf_1166.fifo_rd_block = 0;
    assign fifo_intf_1166.fifo_wr_block = 0;
    assign fifo_intf_1166.finish = finish;
    csv_file_dump fifo_csv_dumper_1166;
    csv_file_dump cstatus_csv_dumper_1166;
    df_fifo_monitor fifo_monitor_1166;
    df_fifo_intf fifo_intf_1167(clock,reset);
    assign fifo_intf_1167.rd_en = AESL_inst_myproject.layer2_out_1166_U.if_read & AESL_inst_myproject.layer2_out_1166_U.if_empty_n;
    assign fifo_intf_1167.wr_en = AESL_inst_myproject.layer2_out_1166_U.if_write & AESL_inst_myproject.layer2_out_1166_U.if_full_n;
    assign fifo_intf_1167.fifo_rd_block = 0;
    assign fifo_intf_1167.fifo_wr_block = 0;
    assign fifo_intf_1167.finish = finish;
    csv_file_dump fifo_csv_dumper_1167;
    csv_file_dump cstatus_csv_dumper_1167;
    df_fifo_monitor fifo_monitor_1167;
    df_fifo_intf fifo_intf_1168(clock,reset);
    assign fifo_intf_1168.rd_en = AESL_inst_myproject.layer2_out_1167_U.if_read & AESL_inst_myproject.layer2_out_1167_U.if_empty_n;
    assign fifo_intf_1168.wr_en = AESL_inst_myproject.layer2_out_1167_U.if_write & AESL_inst_myproject.layer2_out_1167_U.if_full_n;
    assign fifo_intf_1168.fifo_rd_block = 0;
    assign fifo_intf_1168.fifo_wr_block = 0;
    assign fifo_intf_1168.finish = finish;
    csv_file_dump fifo_csv_dumper_1168;
    csv_file_dump cstatus_csv_dumper_1168;
    df_fifo_monitor fifo_monitor_1168;
    df_fifo_intf fifo_intf_1169(clock,reset);
    assign fifo_intf_1169.rd_en = AESL_inst_myproject.layer2_out_1168_U.if_read & AESL_inst_myproject.layer2_out_1168_U.if_empty_n;
    assign fifo_intf_1169.wr_en = AESL_inst_myproject.layer2_out_1168_U.if_write & AESL_inst_myproject.layer2_out_1168_U.if_full_n;
    assign fifo_intf_1169.fifo_rd_block = 0;
    assign fifo_intf_1169.fifo_wr_block = 0;
    assign fifo_intf_1169.finish = finish;
    csv_file_dump fifo_csv_dumper_1169;
    csv_file_dump cstatus_csv_dumper_1169;
    df_fifo_monitor fifo_monitor_1169;
    df_fifo_intf fifo_intf_1170(clock,reset);
    assign fifo_intf_1170.rd_en = AESL_inst_myproject.layer2_out_1169_U.if_read & AESL_inst_myproject.layer2_out_1169_U.if_empty_n;
    assign fifo_intf_1170.wr_en = AESL_inst_myproject.layer2_out_1169_U.if_write & AESL_inst_myproject.layer2_out_1169_U.if_full_n;
    assign fifo_intf_1170.fifo_rd_block = 0;
    assign fifo_intf_1170.fifo_wr_block = 0;
    assign fifo_intf_1170.finish = finish;
    csv_file_dump fifo_csv_dumper_1170;
    csv_file_dump cstatus_csv_dumper_1170;
    df_fifo_monitor fifo_monitor_1170;
    df_fifo_intf fifo_intf_1171(clock,reset);
    assign fifo_intf_1171.rd_en = AESL_inst_myproject.layer2_out_1170_U.if_read & AESL_inst_myproject.layer2_out_1170_U.if_empty_n;
    assign fifo_intf_1171.wr_en = AESL_inst_myproject.layer2_out_1170_U.if_write & AESL_inst_myproject.layer2_out_1170_U.if_full_n;
    assign fifo_intf_1171.fifo_rd_block = 0;
    assign fifo_intf_1171.fifo_wr_block = 0;
    assign fifo_intf_1171.finish = finish;
    csv_file_dump fifo_csv_dumper_1171;
    csv_file_dump cstatus_csv_dumper_1171;
    df_fifo_monitor fifo_monitor_1171;
    df_fifo_intf fifo_intf_1172(clock,reset);
    assign fifo_intf_1172.rd_en = AESL_inst_myproject.layer2_out_1171_U.if_read & AESL_inst_myproject.layer2_out_1171_U.if_empty_n;
    assign fifo_intf_1172.wr_en = AESL_inst_myproject.layer2_out_1171_U.if_write & AESL_inst_myproject.layer2_out_1171_U.if_full_n;
    assign fifo_intf_1172.fifo_rd_block = 0;
    assign fifo_intf_1172.fifo_wr_block = 0;
    assign fifo_intf_1172.finish = finish;
    csv_file_dump fifo_csv_dumper_1172;
    csv_file_dump cstatus_csv_dumper_1172;
    df_fifo_monitor fifo_monitor_1172;
    df_fifo_intf fifo_intf_1173(clock,reset);
    assign fifo_intf_1173.rd_en = AESL_inst_myproject.layer2_out_1172_U.if_read & AESL_inst_myproject.layer2_out_1172_U.if_empty_n;
    assign fifo_intf_1173.wr_en = AESL_inst_myproject.layer2_out_1172_U.if_write & AESL_inst_myproject.layer2_out_1172_U.if_full_n;
    assign fifo_intf_1173.fifo_rd_block = 0;
    assign fifo_intf_1173.fifo_wr_block = 0;
    assign fifo_intf_1173.finish = finish;
    csv_file_dump fifo_csv_dumper_1173;
    csv_file_dump cstatus_csv_dumper_1173;
    df_fifo_monitor fifo_monitor_1173;
    df_fifo_intf fifo_intf_1174(clock,reset);
    assign fifo_intf_1174.rd_en = AESL_inst_myproject.layer2_out_1173_U.if_read & AESL_inst_myproject.layer2_out_1173_U.if_empty_n;
    assign fifo_intf_1174.wr_en = AESL_inst_myproject.layer2_out_1173_U.if_write & AESL_inst_myproject.layer2_out_1173_U.if_full_n;
    assign fifo_intf_1174.fifo_rd_block = 0;
    assign fifo_intf_1174.fifo_wr_block = 0;
    assign fifo_intf_1174.finish = finish;
    csv_file_dump fifo_csv_dumper_1174;
    csv_file_dump cstatus_csv_dumper_1174;
    df_fifo_monitor fifo_monitor_1174;
    df_fifo_intf fifo_intf_1175(clock,reset);
    assign fifo_intf_1175.rd_en = AESL_inst_myproject.layer2_out_1174_U.if_read & AESL_inst_myproject.layer2_out_1174_U.if_empty_n;
    assign fifo_intf_1175.wr_en = AESL_inst_myproject.layer2_out_1174_U.if_write & AESL_inst_myproject.layer2_out_1174_U.if_full_n;
    assign fifo_intf_1175.fifo_rd_block = 0;
    assign fifo_intf_1175.fifo_wr_block = 0;
    assign fifo_intf_1175.finish = finish;
    csv_file_dump fifo_csv_dumper_1175;
    csv_file_dump cstatus_csv_dumper_1175;
    df_fifo_monitor fifo_monitor_1175;
    df_fifo_intf fifo_intf_1176(clock,reset);
    assign fifo_intf_1176.rd_en = AESL_inst_myproject.layer2_out_1175_U.if_read & AESL_inst_myproject.layer2_out_1175_U.if_empty_n;
    assign fifo_intf_1176.wr_en = AESL_inst_myproject.layer2_out_1175_U.if_write & AESL_inst_myproject.layer2_out_1175_U.if_full_n;
    assign fifo_intf_1176.fifo_rd_block = 0;
    assign fifo_intf_1176.fifo_wr_block = 0;
    assign fifo_intf_1176.finish = finish;
    csv_file_dump fifo_csv_dumper_1176;
    csv_file_dump cstatus_csv_dumper_1176;
    df_fifo_monitor fifo_monitor_1176;
    df_fifo_intf fifo_intf_1177(clock,reset);
    assign fifo_intf_1177.rd_en = AESL_inst_myproject.layer2_out_1176_U.if_read & AESL_inst_myproject.layer2_out_1176_U.if_empty_n;
    assign fifo_intf_1177.wr_en = AESL_inst_myproject.layer2_out_1176_U.if_write & AESL_inst_myproject.layer2_out_1176_U.if_full_n;
    assign fifo_intf_1177.fifo_rd_block = 0;
    assign fifo_intf_1177.fifo_wr_block = 0;
    assign fifo_intf_1177.finish = finish;
    csv_file_dump fifo_csv_dumper_1177;
    csv_file_dump cstatus_csv_dumper_1177;
    df_fifo_monitor fifo_monitor_1177;
    df_fifo_intf fifo_intf_1178(clock,reset);
    assign fifo_intf_1178.rd_en = AESL_inst_myproject.layer2_out_1177_U.if_read & AESL_inst_myproject.layer2_out_1177_U.if_empty_n;
    assign fifo_intf_1178.wr_en = AESL_inst_myproject.layer2_out_1177_U.if_write & AESL_inst_myproject.layer2_out_1177_U.if_full_n;
    assign fifo_intf_1178.fifo_rd_block = 0;
    assign fifo_intf_1178.fifo_wr_block = 0;
    assign fifo_intf_1178.finish = finish;
    csv_file_dump fifo_csv_dumper_1178;
    csv_file_dump cstatus_csv_dumper_1178;
    df_fifo_monitor fifo_monitor_1178;
    df_fifo_intf fifo_intf_1179(clock,reset);
    assign fifo_intf_1179.rd_en = AESL_inst_myproject.layer2_out_1178_U.if_read & AESL_inst_myproject.layer2_out_1178_U.if_empty_n;
    assign fifo_intf_1179.wr_en = AESL_inst_myproject.layer2_out_1178_U.if_write & AESL_inst_myproject.layer2_out_1178_U.if_full_n;
    assign fifo_intf_1179.fifo_rd_block = 0;
    assign fifo_intf_1179.fifo_wr_block = 0;
    assign fifo_intf_1179.finish = finish;
    csv_file_dump fifo_csv_dumper_1179;
    csv_file_dump cstatus_csv_dumper_1179;
    df_fifo_monitor fifo_monitor_1179;
    df_fifo_intf fifo_intf_1180(clock,reset);
    assign fifo_intf_1180.rd_en = AESL_inst_myproject.layer2_out_1179_U.if_read & AESL_inst_myproject.layer2_out_1179_U.if_empty_n;
    assign fifo_intf_1180.wr_en = AESL_inst_myproject.layer2_out_1179_U.if_write & AESL_inst_myproject.layer2_out_1179_U.if_full_n;
    assign fifo_intf_1180.fifo_rd_block = 0;
    assign fifo_intf_1180.fifo_wr_block = 0;
    assign fifo_intf_1180.finish = finish;
    csv_file_dump fifo_csv_dumper_1180;
    csv_file_dump cstatus_csv_dumper_1180;
    df_fifo_monitor fifo_monitor_1180;
    df_fifo_intf fifo_intf_1181(clock,reset);
    assign fifo_intf_1181.rd_en = AESL_inst_myproject.layer2_out_1180_U.if_read & AESL_inst_myproject.layer2_out_1180_U.if_empty_n;
    assign fifo_intf_1181.wr_en = AESL_inst_myproject.layer2_out_1180_U.if_write & AESL_inst_myproject.layer2_out_1180_U.if_full_n;
    assign fifo_intf_1181.fifo_rd_block = 0;
    assign fifo_intf_1181.fifo_wr_block = 0;
    assign fifo_intf_1181.finish = finish;
    csv_file_dump fifo_csv_dumper_1181;
    csv_file_dump cstatus_csv_dumper_1181;
    df_fifo_monitor fifo_monitor_1181;
    df_fifo_intf fifo_intf_1182(clock,reset);
    assign fifo_intf_1182.rd_en = AESL_inst_myproject.layer2_out_1181_U.if_read & AESL_inst_myproject.layer2_out_1181_U.if_empty_n;
    assign fifo_intf_1182.wr_en = AESL_inst_myproject.layer2_out_1181_U.if_write & AESL_inst_myproject.layer2_out_1181_U.if_full_n;
    assign fifo_intf_1182.fifo_rd_block = 0;
    assign fifo_intf_1182.fifo_wr_block = 0;
    assign fifo_intf_1182.finish = finish;
    csv_file_dump fifo_csv_dumper_1182;
    csv_file_dump cstatus_csv_dumper_1182;
    df_fifo_monitor fifo_monitor_1182;
    df_fifo_intf fifo_intf_1183(clock,reset);
    assign fifo_intf_1183.rd_en = AESL_inst_myproject.layer2_out_1182_U.if_read & AESL_inst_myproject.layer2_out_1182_U.if_empty_n;
    assign fifo_intf_1183.wr_en = AESL_inst_myproject.layer2_out_1182_U.if_write & AESL_inst_myproject.layer2_out_1182_U.if_full_n;
    assign fifo_intf_1183.fifo_rd_block = 0;
    assign fifo_intf_1183.fifo_wr_block = 0;
    assign fifo_intf_1183.finish = finish;
    csv_file_dump fifo_csv_dumper_1183;
    csv_file_dump cstatus_csv_dumper_1183;
    df_fifo_monitor fifo_monitor_1183;
    df_fifo_intf fifo_intf_1184(clock,reset);
    assign fifo_intf_1184.rd_en = AESL_inst_myproject.layer2_out_1183_U.if_read & AESL_inst_myproject.layer2_out_1183_U.if_empty_n;
    assign fifo_intf_1184.wr_en = AESL_inst_myproject.layer2_out_1183_U.if_write & AESL_inst_myproject.layer2_out_1183_U.if_full_n;
    assign fifo_intf_1184.fifo_rd_block = 0;
    assign fifo_intf_1184.fifo_wr_block = 0;
    assign fifo_intf_1184.finish = finish;
    csv_file_dump fifo_csv_dumper_1184;
    csv_file_dump cstatus_csv_dumper_1184;
    df_fifo_monitor fifo_monitor_1184;
    df_fifo_intf fifo_intf_1185(clock,reset);
    assign fifo_intf_1185.rd_en = AESL_inst_myproject.layer2_out_1184_U.if_read & AESL_inst_myproject.layer2_out_1184_U.if_empty_n;
    assign fifo_intf_1185.wr_en = AESL_inst_myproject.layer2_out_1184_U.if_write & AESL_inst_myproject.layer2_out_1184_U.if_full_n;
    assign fifo_intf_1185.fifo_rd_block = 0;
    assign fifo_intf_1185.fifo_wr_block = 0;
    assign fifo_intf_1185.finish = finish;
    csv_file_dump fifo_csv_dumper_1185;
    csv_file_dump cstatus_csv_dumper_1185;
    df_fifo_monitor fifo_monitor_1185;
    df_fifo_intf fifo_intf_1186(clock,reset);
    assign fifo_intf_1186.rd_en = AESL_inst_myproject.layer2_out_1185_U.if_read & AESL_inst_myproject.layer2_out_1185_U.if_empty_n;
    assign fifo_intf_1186.wr_en = AESL_inst_myproject.layer2_out_1185_U.if_write & AESL_inst_myproject.layer2_out_1185_U.if_full_n;
    assign fifo_intf_1186.fifo_rd_block = 0;
    assign fifo_intf_1186.fifo_wr_block = 0;
    assign fifo_intf_1186.finish = finish;
    csv_file_dump fifo_csv_dumper_1186;
    csv_file_dump cstatus_csv_dumper_1186;
    df_fifo_monitor fifo_monitor_1186;
    df_fifo_intf fifo_intf_1187(clock,reset);
    assign fifo_intf_1187.rd_en = AESL_inst_myproject.layer2_out_1186_U.if_read & AESL_inst_myproject.layer2_out_1186_U.if_empty_n;
    assign fifo_intf_1187.wr_en = AESL_inst_myproject.layer2_out_1186_U.if_write & AESL_inst_myproject.layer2_out_1186_U.if_full_n;
    assign fifo_intf_1187.fifo_rd_block = 0;
    assign fifo_intf_1187.fifo_wr_block = 0;
    assign fifo_intf_1187.finish = finish;
    csv_file_dump fifo_csv_dumper_1187;
    csv_file_dump cstatus_csv_dumper_1187;
    df_fifo_monitor fifo_monitor_1187;
    df_fifo_intf fifo_intf_1188(clock,reset);
    assign fifo_intf_1188.rd_en = AESL_inst_myproject.layer2_out_1187_U.if_read & AESL_inst_myproject.layer2_out_1187_U.if_empty_n;
    assign fifo_intf_1188.wr_en = AESL_inst_myproject.layer2_out_1187_U.if_write & AESL_inst_myproject.layer2_out_1187_U.if_full_n;
    assign fifo_intf_1188.fifo_rd_block = 0;
    assign fifo_intf_1188.fifo_wr_block = 0;
    assign fifo_intf_1188.finish = finish;
    csv_file_dump fifo_csv_dumper_1188;
    csv_file_dump cstatus_csv_dumper_1188;
    df_fifo_monitor fifo_monitor_1188;
    df_fifo_intf fifo_intf_1189(clock,reset);
    assign fifo_intf_1189.rd_en = AESL_inst_myproject.layer2_out_1188_U.if_read & AESL_inst_myproject.layer2_out_1188_U.if_empty_n;
    assign fifo_intf_1189.wr_en = AESL_inst_myproject.layer2_out_1188_U.if_write & AESL_inst_myproject.layer2_out_1188_U.if_full_n;
    assign fifo_intf_1189.fifo_rd_block = 0;
    assign fifo_intf_1189.fifo_wr_block = 0;
    assign fifo_intf_1189.finish = finish;
    csv_file_dump fifo_csv_dumper_1189;
    csv_file_dump cstatus_csv_dumper_1189;
    df_fifo_monitor fifo_monitor_1189;
    df_fifo_intf fifo_intf_1190(clock,reset);
    assign fifo_intf_1190.rd_en = AESL_inst_myproject.layer2_out_1189_U.if_read & AESL_inst_myproject.layer2_out_1189_U.if_empty_n;
    assign fifo_intf_1190.wr_en = AESL_inst_myproject.layer2_out_1189_U.if_write & AESL_inst_myproject.layer2_out_1189_U.if_full_n;
    assign fifo_intf_1190.fifo_rd_block = 0;
    assign fifo_intf_1190.fifo_wr_block = 0;
    assign fifo_intf_1190.finish = finish;
    csv_file_dump fifo_csv_dumper_1190;
    csv_file_dump cstatus_csv_dumper_1190;
    df_fifo_monitor fifo_monitor_1190;
    df_fifo_intf fifo_intf_1191(clock,reset);
    assign fifo_intf_1191.rd_en = AESL_inst_myproject.layer2_out_1190_U.if_read & AESL_inst_myproject.layer2_out_1190_U.if_empty_n;
    assign fifo_intf_1191.wr_en = AESL_inst_myproject.layer2_out_1190_U.if_write & AESL_inst_myproject.layer2_out_1190_U.if_full_n;
    assign fifo_intf_1191.fifo_rd_block = 0;
    assign fifo_intf_1191.fifo_wr_block = 0;
    assign fifo_intf_1191.finish = finish;
    csv_file_dump fifo_csv_dumper_1191;
    csv_file_dump cstatus_csv_dumper_1191;
    df_fifo_monitor fifo_monitor_1191;
    df_fifo_intf fifo_intf_1192(clock,reset);
    assign fifo_intf_1192.rd_en = AESL_inst_myproject.layer2_out_1191_U.if_read & AESL_inst_myproject.layer2_out_1191_U.if_empty_n;
    assign fifo_intf_1192.wr_en = AESL_inst_myproject.layer2_out_1191_U.if_write & AESL_inst_myproject.layer2_out_1191_U.if_full_n;
    assign fifo_intf_1192.fifo_rd_block = 0;
    assign fifo_intf_1192.fifo_wr_block = 0;
    assign fifo_intf_1192.finish = finish;
    csv_file_dump fifo_csv_dumper_1192;
    csv_file_dump cstatus_csv_dumper_1192;
    df_fifo_monitor fifo_monitor_1192;
    df_fifo_intf fifo_intf_1193(clock,reset);
    assign fifo_intf_1193.rd_en = AESL_inst_myproject.layer2_out_1192_U.if_read & AESL_inst_myproject.layer2_out_1192_U.if_empty_n;
    assign fifo_intf_1193.wr_en = AESL_inst_myproject.layer2_out_1192_U.if_write & AESL_inst_myproject.layer2_out_1192_U.if_full_n;
    assign fifo_intf_1193.fifo_rd_block = 0;
    assign fifo_intf_1193.fifo_wr_block = 0;
    assign fifo_intf_1193.finish = finish;
    csv_file_dump fifo_csv_dumper_1193;
    csv_file_dump cstatus_csv_dumper_1193;
    df_fifo_monitor fifo_monitor_1193;
    df_fifo_intf fifo_intf_1194(clock,reset);
    assign fifo_intf_1194.rd_en = AESL_inst_myproject.layer2_out_1193_U.if_read & AESL_inst_myproject.layer2_out_1193_U.if_empty_n;
    assign fifo_intf_1194.wr_en = AESL_inst_myproject.layer2_out_1193_U.if_write & AESL_inst_myproject.layer2_out_1193_U.if_full_n;
    assign fifo_intf_1194.fifo_rd_block = 0;
    assign fifo_intf_1194.fifo_wr_block = 0;
    assign fifo_intf_1194.finish = finish;
    csv_file_dump fifo_csv_dumper_1194;
    csv_file_dump cstatus_csv_dumper_1194;
    df_fifo_monitor fifo_monitor_1194;
    df_fifo_intf fifo_intf_1195(clock,reset);
    assign fifo_intf_1195.rd_en = AESL_inst_myproject.layer2_out_1194_U.if_read & AESL_inst_myproject.layer2_out_1194_U.if_empty_n;
    assign fifo_intf_1195.wr_en = AESL_inst_myproject.layer2_out_1194_U.if_write & AESL_inst_myproject.layer2_out_1194_U.if_full_n;
    assign fifo_intf_1195.fifo_rd_block = 0;
    assign fifo_intf_1195.fifo_wr_block = 0;
    assign fifo_intf_1195.finish = finish;
    csv_file_dump fifo_csv_dumper_1195;
    csv_file_dump cstatus_csv_dumper_1195;
    df_fifo_monitor fifo_monitor_1195;
    df_fifo_intf fifo_intf_1196(clock,reset);
    assign fifo_intf_1196.rd_en = AESL_inst_myproject.layer2_out_1195_U.if_read & AESL_inst_myproject.layer2_out_1195_U.if_empty_n;
    assign fifo_intf_1196.wr_en = AESL_inst_myproject.layer2_out_1195_U.if_write & AESL_inst_myproject.layer2_out_1195_U.if_full_n;
    assign fifo_intf_1196.fifo_rd_block = 0;
    assign fifo_intf_1196.fifo_wr_block = 0;
    assign fifo_intf_1196.finish = finish;
    csv_file_dump fifo_csv_dumper_1196;
    csv_file_dump cstatus_csv_dumper_1196;
    df_fifo_monitor fifo_monitor_1196;
    df_fifo_intf fifo_intf_1197(clock,reset);
    assign fifo_intf_1197.rd_en = AESL_inst_myproject.layer2_out_1196_U.if_read & AESL_inst_myproject.layer2_out_1196_U.if_empty_n;
    assign fifo_intf_1197.wr_en = AESL_inst_myproject.layer2_out_1196_U.if_write & AESL_inst_myproject.layer2_out_1196_U.if_full_n;
    assign fifo_intf_1197.fifo_rd_block = 0;
    assign fifo_intf_1197.fifo_wr_block = 0;
    assign fifo_intf_1197.finish = finish;
    csv_file_dump fifo_csv_dumper_1197;
    csv_file_dump cstatus_csv_dumper_1197;
    df_fifo_monitor fifo_monitor_1197;
    df_fifo_intf fifo_intf_1198(clock,reset);
    assign fifo_intf_1198.rd_en = AESL_inst_myproject.layer2_out_1197_U.if_read & AESL_inst_myproject.layer2_out_1197_U.if_empty_n;
    assign fifo_intf_1198.wr_en = AESL_inst_myproject.layer2_out_1197_U.if_write & AESL_inst_myproject.layer2_out_1197_U.if_full_n;
    assign fifo_intf_1198.fifo_rd_block = 0;
    assign fifo_intf_1198.fifo_wr_block = 0;
    assign fifo_intf_1198.finish = finish;
    csv_file_dump fifo_csv_dumper_1198;
    csv_file_dump cstatus_csv_dumper_1198;
    df_fifo_monitor fifo_monitor_1198;
    df_fifo_intf fifo_intf_1199(clock,reset);
    assign fifo_intf_1199.rd_en = AESL_inst_myproject.layer2_out_1198_U.if_read & AESL_inst_myproject.layer2_out_1198_U.if_empty_n;
    assign fifo_intf_1199.wr_en = AESL_inst_myproject.layer2_out_1198_U.if_write & AESL_inst_myproject.layer2_out_1198_U.if_full_n;
    assign fifo_intf_1199.fifo_rd_block = 0;
    assign fifo_intf_1199.fifo_wr_block = 0;
    assign fifo_intf_1199.finish = finish;
    csv_file_dump fifo_csv_dumper_1199;
    csv_file_dump cstatus_csv_dumper_1199;
    df_fifo_monitor fifo_monitor_1199;
    df_fifo_intf fifo_intf_1200(clock,reset);
    assign fifo_intf_1200.rd_en = AESL_inst_myproject.layer2_out_1199_U.if_read & AESL_inst_myproject.layer2_out_1199_U.if_empty_n;
    assign fifo_intf_1200.wr_en = AESL_inst_myproject.layer2_out_1199_U.if_write & AESL_inst_myproject.layer2_out_1199_U.if_full_n;
    assign fifo_intf_1200.fifo_rd_block = 0;
    assign fifo_intf_1200.fifo_wr_block = 0;
    assign fifo_intf_1200.finish = finish;
    csv_file_dump fifo_csv_dumper_1200;
    csv_file_dump cstatus_csv_dumper_1200;
    df_fifo_monitor fifo_monitor_1200;
    df_fifo_intf fifo_intf_1201(clock,reset);
    assign fifo_intf_1201.rd_en = AESL_inst_myproject.layer2_out_1200_U.if_read & AESL_inst_myproject.layer2_out_1200_U.if_empty_n;
    assign fifo_intf_1201.wr_en = AESL_inst_myproject.layer2_out_1200_U.if_write & AESL_inst_myproject.layer2_out_1200_U.if_full_n;
    assign fifo_intf_1201.fifo_rd_block = 0;
    assign fifo_intf_1201.fifo_wr_block = 0;
    assign fifo_intf_1201.finish = finish;
    csv_file_dump fifo_csv_dumper_1201;
    csv_file_dump cstatus_csv_dumper_1201;
    df_fifo_monitor fifo_monitor_1201;
    df_fifo_intf fifo_intf_1202(clock,reset);
    assign fifo_intf_1202.rd_en = AESL_inst_myproject.layer2_out_1201_U.if_read & AESL_inst_myproject.layer2_out_1201_U.if_empty_n;
    assign fifo_intf_1202.wr_en = AESL_inst_myproject.layer2_out_1201_U.if_write & AESL_inst_myproject.layer2_out_1201_U.if_full_n;
    assign fifo_intf_1202.fifo_rd_block = 0;
    assign fifo_intf_1202.fifo_wr_block = 0;
    assign fifo_intf_1202.finish = finish;
    csv_file_dump fifo_csv_dumper_1202;
    csv_file_dump cstatus_csv_dumper_1202;
    df_fifo_monitor fifo_monitor_1202;
    df_fifo_intf fifo_intf_1203(clock,reset);
    assign fifo_intf_1203.rd_en = AESL_inst_myproject.layer2_out_1202_U.if_read & AESL_inst_myproject.layer2_out_1202_U.if_empty_n;
    assign fifo_intf_1203.wr_en = AESL_inst_myproject.layer2_out_1202_U.if_write & AESL_inst_myproject.layer2_out_1202_U.if_full_n;
    assign fifo_intf_1203.fifo_rd_block = 0;
    assign fifo_intf_1203.fifo_wr_block = 0;
    assign fifo_intf_1203.finish = finish;
    csv_file_dump fifo_csv_dumper_1203;
    csv_file_dump cstatus_csv_dumper_1203;
    df_fifo_monitor fifo_monitor_1203;
    df_fifo_intf fifo_intf_1204(clock,reset);
    assign fifo_intf_1204.rd_en = AESL_inst_myproject.layer2_out_1203_U.if_read & AESL_inst_myproject.layer2_out_1203_U.if_empty_n;
    assign fifo_intf_1204.wr_en = AESL_inst_myproject.layer2_out_1203_U.if_write & AESL_inst_myproject.layer2_out_1203_U.if_full_n;
    assign fifo_intf_1204.fifo_rd_block = 0;
    assign fifo_intf_1204.fifo_wr_block = 0;
    assign fifo_intf_1204.finish = finish;
    csv_file_dump fifo_csv_dumper_1204;
    csv_file_dump cstatus_csv_dumper_1204;
    df_fifo_monitor fifo_monitor_1204;
    df_fifo_intf fifo_intf_1205(clock,reset);
    assign fifo_intf_1205.rd_en = AESL_inst_myproject.layer2_out_1204_U.if_read & AESL_inst_myproject.layer2_out_1204_U.if_empty_n;
    assign fifo_intf_1205.wr_en = AESL_inst_myproject.layer2_out_1204_U.if_write & AESL_inst_myproject.layer2_out_1204_U.if_full_n;
    assign fifo_intf_1205.fifo_rd_block = 0;
    assign fifo_intf_1205.fifo_wr_block = 0;
    assign fifo_intf_1205.finish = finish;
    csv_file_dump fifo_csv_dumper_1205;
    csv_file_dump cstatus_csv_dumper_1205;
    df_fifo_monitor fifo_monitor_1205;
    df_fifo_intf fifo_intf_1206(clock,reset);
    assign fifo_intf_1206.rd_en = AESL_inst_myproject.layer2_out_1205_U.if_read & AESL_inst_myproject.layer2_out_1205_U.if_empty_n;
    assign fifo_intf_1206.wr_en = AESL_inst_myproject.layer2_out_1205_U.if_write & AESL_inst_myproject.layer2_out_1205_U.if_full_n;
    assign fifo_intf_1206.fifo_rd_block = 0;
    assign fifo_intf_1206.fifo_wr_block = 0;
    assign fifo_intf_1206.finish = finish;
    csv_file_dump fifo_csv_dumper_1206;
    csv_file_dump cstatus_csv_dumper_1206;
    df_fifo_monitor fifo_monitor_1206;
    df_fifo_intf fifo_intf_1207(clock,reset);
    assign fifo_intf_1207.rd_en = AESL_inst_myproject.layer2_out_1206_U.if_read & AESL_inst_myproject.layer2_out_1206_U.if_empty_n;
    assign fifo_intf_1207.wr_en = AESL_inst_myproject.layer2_out_1206_U.if_write & AESL_inst_myproject.layer2_out_1206_U.if_full_n;
    assign fifo_intf_1207.fifo_rd_block = 0;
    assign fifo_intf_1207.fifo_wr_block = 0;
    assign fifo_intf_1207.finish = finish;
    csv_file_dump fifo_csv_dumper_1207;
    csv_file_dump cstatus_csv_dumper_1207;
    df_fifo_monitor fifo_monitor_1207;
    df_fifo_intf fifo_intf_1208(clock,reset);
    assign fifo_intf_1208.rd_en = AESL_inst_myproject.layer2_out_1207_U.if_read & AESL_inst_myproject.layer2_out_1207_U.if_empty_n;
    assign fifo_intf_1208.wr_en = AESL_inst_myproject.layer2_out_1207_U.if_write & AESL_inst_myproject.layer2_out_1207_U.if_full_n;
    assign fifo_intf_1208.fifo_rd_block = 0;
    assign fifo_intf_1208.fifo_wr_block = 0;
    assign fifo_intf_1208.finish = finish;
    csv_file_dump fifo_csv_dumper_1208;
    csv_file_dump cstatus_csv_dumper_1208;
    df_fifo_monitor fifo_monitor_1208;
    df_fifo_intf fifo_intf_1209(clock,reset);
    assign fifo_intf_1209.rd_en = AESL_inst_myproject.layer2_out_1208_U.if_read & AESL_inst_myproject.layer2_out_1208_U.if_empty_n;
    assign fifo_intf_1209.wr_en = AESL_inst_myproject.layer2_out_1208_U.if_write & AESL_inst_myproject.layer2_out_1208_U.if_full_n;
    assign fifo_intf_1209.fifo_rd_block = 0;
    assign fifo_intf_1209.fifo_wr_block = 0;
    assign fifo_intf_1209.finish = finish;
    csv_file_dump fifo_csv_dumper_1209;
    csv_file_dump cstatus_csv_dumper_1209;
    df_fifo_monitor fifo_monitor_1209;
    df_fifo_intf fifo_intf_1210(clock,reset);
    assign fifo_intf_1210.rd_en = AESL_inst_myproject.layer2_out_1209_U.if_read & AESL_inst_myproject.layer2_out_1209_U.if_empty_n;
    assign fifo_intf_1210.wr_en = AESL_inst_myproject.layer2_out_1209_U.if_write & AESL_inst_myproject.layer2_out_1209_U.if_full_n;
    assign fifo_intf_1210.fifo_rd_block = 0;
    assign fifo_intf_1210.fifo_wr_block = 0;
    assign fifo_intf_1210.finish = finish;
    csv_file_dump fifo_csv_dumper_1210;
    csv_file_dump cstatus_csv_dumper_1210;
    df_fifo_monitor fifo_monitor_1210;
    df_fifo_intf fifo_intf_1211(clock,reset);
    assign fifo_intf_1211.rd_en = AESL_inst_myproject.layer2_out_1210_U.if_read & AESL_inst_myproject.layer2_out_1210_U.if_empty_n;
    assign fifo_intf_1211.wr_en = AESL_inst_myproject.layer2_out_1210_U.if_write & AESL_inst_myproject.layer2_out_1210_U.if_full_n;
    assign fifo_intf_1211.fifo_rd_block = 0;
    assign fifo_intf_1211.fifo_wr_block = 0;
    assign fifo_intf_1211.finish = finish;
    csv_file_dump fifo_csv_dumper_1211;
    csv_file_dump cstatus_csv_dumper_1211;
    df_fifo_monitor fifo_monitor_1211;
    df_fifo_intf fifo_intf_1212(clock,reset);
    assign fifo_intf_1212.rd_en = AESL_inst_myproject.layer2_out_1211_U.if_read & AESL_inst_myproject.layer2_out_1211_U.if_empty_n;
    assign fifo_intf_1212.wr_en = AESL_inst_myproject.layer2_out_1211_U.if_write & AESL_inst_myproject.layer2_out_1211_U.if_full_n;
    assign fifo_intf_1212.fifo_rd_block = 0;
    assign fifo_intf_1212.fifo_wr_block = 0;
    assign fifo_intf_1212.finish = finish;
    csv_file_dump fifo_csv_dumper_1212;
    csv_file_dump cstatus_csv_dumper_1212;
    df_fifo_monitor fifo_monitor_1212;
    df_fifo_intf fifo_intf_1213(clock,reset);
    assign fifo_intf_1213.rd_en = AESL_inst_myproject.layer2_out_1212_U.if_read & AESL_inst_myproject.layer2_out_1212_U.if_empty_n;
    assign fifo_intf_1213.wr_en = AESL_inst_myproject.layer2_out_1212_U.if_write & AESL_inst_myproject.layer2_out_1212_U.if_full_n;
    assign fifo_intf_1213.fifo_rd_block = 0;
    assign fifo_intf_1213.fifo_wr_block = 0;
    assign fifo_intf_1213.finish = finish;
    csv_file_dump fifo_csv_dumper_1213;
    csv_file_dump cstatus_csv_dumper_1213;
    df_fifo_monitor fifo_monitor_1213;
    df_fifo_intf fifo_intf_1214(clock,reset);
    assign fifo_intf_1214.rd_en = AESL_inst_myproject.layer2_out_1213_U.if_read & AESL_inst_myproject.layer2_out_1213_U.if_empty_n;
    assign fifo_intf_1214.wr_en = AESL_inst_myproject.layer2_out_1213_U.if_write & AESL_inst_myproject.layer2_out_1213_U.if_full_n;
    assign fifo_intf_1214.fifo_rd_block = 0;
    assign fifo_intf_1214.fifo_wr_block = 0;
    assign fifo_intf_1214.finish = finish;
    csv_file_dump fifo_csv_dumper_1214;
    csv_file_dump cstatus_csv_dumper_1214;
    df_fifo_monitor fifo_monitor_1214;
    df_fifo_intf fifo_intf_1215(clock,reset);
    assign fifo_intf_1215.rd_en = AESL_inst_myproject.layer2_out_1214_U.if_read & AESL_inst_myproject.layer2_out_1214_U.if_empty_n;
    assign fifo_intf_1215.wr_en = AESL_inst_myproject.layer2_out_1214_U.if_write & AESL_inst_myproject.layer2_out_1214_U.if_full_n;
    assign fifo_intf_1215.fifo_rd_block = 0;
    assign fifo_intf_1215.fifo_wr_block = 0;
    assign fifo_intf_1215.finish = finish;
    csv_file_dump fifo_csv_dumper_1215;
    csv_file_dump cstatus_csv_dumper_1215;
    df_fifo_monitor fifo_monitor_1215;
    df_fifo_intf fifo_intf_1216(clock,reset);
    assign fifo_intf_1216.rd_en = AESL_inst_myproject.layer2_out_1215_U.if_read & AESL_inst_myproject.layer2_out_1215_U.if_empty_n;
    assign fifo_intf_1216.wr_en = AESL_inst_myproject.layer2_out_1215_U.if_write & AESL_inst_myproject.layer2_out_1215_U.if_full_n;
    assign fifo_intf_1216.fifo_rd_block = 0;
    assign fifo_intf_1216.fifo_wr_block = 0;
    assign fifo_intf_1216.finish = finish;
    csv_file_dump fifo_csv_dumper_1216;
    csv_file_dump cstatus_csv_dumper_1216;
    df_fifo_monitor fifo_monitor_1216;
    df_fifo_intf fifo_intf_1217(clock,reset);
    assign fifo_intf_1217.rd_en = AESL_inst_myproject.layer2_out_1216_U.if_read & AESL_inst_myproject.layer2_out_1216_U.if_empty_n;
    assign fifo_intf_1217.wr_en = AESL_inst_myproject.layer2_out_1216_U.if_write & AESL_inst_myproject.layer2_out_1216_U.if_full_n;
    assign fifo_intf_1217.fifo_rd_block = 0;
    assign fifo_intf_1217.fifo_wr_block = 0;
    assign fifo_intf_1217.finish = finish;
    csv_file_dump fifo_csv_dumper_1217;
    csv_file_dump cstatus_csv_dumper_1217;
    df_fifo_monitor fifo_monitor_1217;
    df_fifo_intf fifo_intf_1218(clock,reset);
    assign fifo_intf_1218.rd_en = AESL_inst_myproject.layer2_out_1217_U.if_read & AESL_inst_myproject.layer2_out_1217_U.if_empty_n;
    assign fifo_intf_1218.wr_en = AESL_inst_myproject.layer2_out_1217_U.if_write & AESL_inst_myproject.layer2_out_1217_U.if_full_n;
    assign fifo_intf_1218.fifo_rd_block = 0;
    assign fifo_intf_1218.fifo_wr_block = 0;
    assign fifo_intf_1218.finish = finish;
    csv_file_dump fifo_csv_dumper_1218;
    csv_file_dump cstatus_csv_dumper_1218;
    df_fifo_monitor fifo_monitor_1218;
    df_fifo_intf fifo_intf_1219(clock,reset);
    assign fifo_intf_1219.rd_en = AESL_inst_myproject.layer2_out_1218_U.if_read & AESL_inst_myproject.layer2_out_1218_U.if_empty_n;
    assign fifo_intf_1219.wr_en = AESL_inst_myproject.layer2_out_1218_U.if_write & AESL_inst_myproject.layer2_out_1218_U.if_full_n;
    assign fifo_intf_1219.fifo_rd_block = 0;
    assign fifo_intf_1219.fifo_wr_block = 0;
    assign fifo_intf_1219.finish = finish;
    csv_file_dump fifo_csv_dumper_1219;
    csv_file_dump cstatus_csv_dumper_1219;
    df_fifo_monitor fifo_monitor_1219;
    df_fifo_intf fifo_intf_1220(clock,reset);
    assign fifo_intf_1220.rd_en = AESL_inst_myproject.layer2_out_1219_U.if_read & AESL_inst_myproject.layer2_out_1219_U.if_empty_n;
    assign fifo_intf_1220.wr_en = AESL_inst_myproject.layer2_out_1219_U.if_write & AESL_inst_myproject.layer2_out_1219_U.if_full_n;
    assign fifo_intf_1220.fifo_rd_block = 0;
    assign fifo_intf_1220.fifo_wr_block = 0;
    assign fifo_intf_1220.finish = finish;
    csv_file_dump fifo_csv_dumper_1220;
    csv_file_dump cstatus_csv_dumper_1220;
    df_fifo_monitor fifo_monitor_1220;
    df_fifo_intf fifo_intf_1221(clock,reset);
    assign fifo_intf_1221.rd_en = AESL_inst_myproject.layer2_out_1220_U.if_read & AESL_inst_myproject.layer2_out_1220_U.if_empty_n;
    assign fifo_intf_1221.wr_en = AESL_inst_myproject.layer2_out_1220_U.if_write & AESL_inst_myproject.layer2_out_1220_U.if_full_n;
    assign fifo_intf_1221.fifo_rd_block = 0;
    assign fifo_intf_1221.fifo_wr_block = 0;
    assign fifo_intf_1221.finish = finish;
    csv_file_dump fifo_csv_dumper_1221;
    csv_file_dump cstatus_csv_dumper_1221;
    df_fifo_monitor fifo_monitor_1221;
    df_fifo_intf fifo_intf_1222(clock,reset);
    assign fifo_intf_1222.rd_en = AESL_inst_myproject.layer2_out_1221_U.if_read & AESL_inst_myproject.layer2_out_1221_U.if_empty_n;
    assign fifo_intf_1222.wr_en = AESL_inst_myproject.layer2_out_1221_U.if_write & AESL_inst_myproject.layer2_out_1221_U.if_full_n;
    assign fifo_intf_1222.fifo_rd_block = 0;
    assign fifo_intf_1222.fifo_wr_block = 0;
    assign fifo_intf_1222.finish = finish;
    csv_file_dump fifo_csv_dumper_1222;
    csv_file_dump cstatus_csv_dumper_1222;
    df_fifo_monitor fifo_monitor_1222;
    df_fifo_intf fifo_intf_1223(clock,reset);
    assign fifo_intf_1223.rd_en = AESL_inst_myproject.layer2_out_1222_U.if_read & AESL_inst_myproject.layer2_out_1222_U.if_empty_n;
    assign fifo_intf_1223.wr_en = AESL_inst_myproject.layer2_out_1222_U.if_write & AESL_inst_myproject.layer2_out_1222_U.if_full_n;
    assign fifo_intf_1223.fifo_rd_block = 0;
    assign fifo_intf_1223.fifo_wr_block = 0;
    assign fifo_intf_1223.finish = finish;
    csv_file_dump fifo_csv_dumper_1223;
    csv_file_dump cstatus_csv_dumper_1223;
    df_fifo_monitor fifo_monitor_1223;
    df_fifo_intf fifo_intf_1224(clock,reset);
    assign fifo_intf_1224.rd_en = AESL_inst_myproject.layer2_out_1223_U.if_read & AESL_inst_myproject.layer2_out_1223_U.if_empty_n;
    assign fifo_intf_1224.wr_en = AESL_inst_myproject.layer2_out_1223_U.if_write & AESL_inst_myproject.layer2_out_1223_U.if_full_n;
    assign fifo_intf_1224.fifo_rd_block = 0;
    assign fifo_intf_1224.fifo_wr_block = 0;
    assign fifo_intf_1224.finish = finish;
    csv_file_dump fifo_csv_dumper_1224;
    csv_file_dump cstatus_csv_dumper_1224;
    df_fifo_monitor fifo_monitor_1224;
    df_fifo_intf fifo_intf_1225(clock,reset);
    assign fifo_intf_1225.rd_en = AESL_inst_myproject.layer2_out_1224_U.if_read & AESL_inst_myproject.layer2_out_1224_U.if_empty_n;
    assign fifo_intf_1225.wr_en = AESL_inst_myproject.layer2_out_1224_U.if_write & AESL_inst_myproject.layer2_out_1224_U.if_full_n;
    assign fifo_intf_1225.fifo_rd_block = 0;
    assign fifo_intf_1225.fifo_wr_block = 0;
    assign fifo_intf_1225.finish = finish;
    csv_file_dump fifo_csv_dumper_1225;
    csv_file_dump cstatus_csv_dumper_1225;
    df_fifo_monitor fifo_monitor_1225;
    df_fifo_intf fifo_intf_1226(clock,reset);
    assign fifo_intf_1226.rd_en = AESL_inst_myproject.layer2_out_1225_U.if_read & AESL_inst_myproject.layer2_out_1225_U.if_empty_n;
    assign fifo_intf_1226.wr_en = AESL_inst_myproject.layer2_out_1225_U.if_write & AESL_inst_myproject.layer2_out_1225_U.if_full_n;
    assign fifo_intf_1226.fifo_rd_block = 0;
    assign fifo_intf_1226.fifo_wr_block = 0;
    assign fifo_intf_1226.finish = finish;
    csv_file_dump fifo_csv_dumper_1226;
    csv_file_dump cstatus_csv_dumper_1226;
    df_fifo_monitor fifo_monitor_1226;
    df_fifo_intf fifo_intf_1227(clock,reset);
    assign fifo_intf_1227.rd_en = AESL_inst_myproject.layer2_out_1226_U.if_read & AESL_inst_myproject.layer2_out_1226_U.if_empty_n;
    assign fifo_intf_1227.wr_en = AESL_inst_myproject.layer2_out_1226_U.if_write & AESL_inst_myproject.layer2_out_1226_U.if_full_n;
    assign fifo_intf_1227.fifo_rd_block = 0;
    assign fifo_intf_1227.fifo_wr_block = 0;
    assign fifo_intf_1227.finish = finish;
    csv_file_dump fifo_csv_dumper_1227;
    csv_file_dump cstatus_csv_dumper_1227;
    df_fifo_monitor fifo_monitor_1227;
    df_fifo_intf fifo_intf_1228(clock,reset);
    assign fifo_intf_1228.rd_en = AESL_inst_myproject.layer2_out_1227_U.if_read & AESL_inst_myproject.layer2_out_1227_U.if_empty_n;
    assign fifo_intf_1228.wr_en = AESL_inst_myproject.layer2_out_1227_U.if_write & AESL_inst_myproject.layer2_out_1227_U.if_full_n;
    assign fifo_intf_1228.fifo_rd_block = 0;
    assign fifo_intf_1228.fifo_wr_block = 0;
    assign fifo_intf_1228.finish = finish;
    csv_file_dump fifo_csv_dumper_1228;
    csv_file_dump cstatus_csv_dumper_1228;
    df_fifo_monitor fifo_monitor_1228;
    df_fifo_intf fifo_intf_1229(clock,reset);
    assign fifo_intf_1229.rd_en = AESL_inst_myproject.layer2_out_1228_U.if_read & AESL_inst_myproject.layer2_out_1228_U.if_empty_n;
    assign fifo_intf_1229.wr_en = AESL_inst_myproject.layer2_out_1228_U.if_write & AESL_inst_myproject.layer2_out_1228_U.if_full_n;
    assign fifo_intf_1229.fifo_rd_block = 0;
    assign fifo_intf_1229.fifo_wr_block = 0;
    assign fifo_intf_1229.finish = finish;
    csv_file_dump fifo_csv_dumper_1229;
    csv_file_dump cstatus_csv_dumper_1229;
    df_fifo_monitor fifo_monitor_1229;
    df_fifo_intf fifo_intf_1230(clock,reset);
    assign fifo_intf_1230.rd_en = AESL_inst_myproject.layer2_out_1229_U.if_read & AESL_inst_myproject.layer2_out_1229_U.if_empty_n;
    assign fifo_intf_1230.wr_en = AESL_inst_myproject.layer2_out_1229_U.if_write & AESL_inst_myproject.layer2_out_1229_U.if_full_n;
    assign fifo_intf_1230.fifo_rd_block = 0;
    assign fifo_intf_1230.fifo_wr_block = 0;
    assign fifo_intf_1230.finish = finish;
    csv_file_dump fifo_csv_dumper_1230;
    csv_file_dump cstatus_csv_dumper_1230;
    df_fifo_monitor fifo_monitor_1230;
    df_fifo_intf fifo_intf_1231(clock,reset);
    assign fifo_intf_1231.rd_en = AESL_inst_myproject.layer2_out_1230_U.if_read & AESL_inst_myproject.layer2_out_1230_U.if_empty_n;
    assign fifo_intf_1231.wr_en = AESL_inst_myproject.layer2_out_1230_U.if_write & AESL_inst_myproject.layer2_out_1230_U.if_full_n;
    assign fifo_intf_1231.fifo_rd_block = 0;
    assign fifo_intf_1231.fifo_wr_block = 0;
    assign fifo_intf_1231.finish = finish;
    csv_file_dump fifo_csv_dumper_1231;
    csv_file_dump cstatus_csv_dumper_1231;
    df_fifo_monitor fifo_monitor_1231;
    df_fifo_intf fifo_intf_1232(clock,reset);
    assign fifo_intf_1232.rd_en = AESL_inst_myproject.layer2_out_1231_U.if_read & AESL_inst_myproject.layer2_out_1231_U.if_empty_n;
    assign fifo_intf_1232.wr_en = AESL_inst_myproject.layer2_out_1231_U.if_write & AESL_inst_myproject.layer2_out_1231_U.if_full_n;
    assign fifo_intf_1232.fifo_rd_block = 0;
    assign fifo_intf_1232.fifo_wr_block = 0;
    assign fifo_intf_1232.finish = finish;
    csv_file_dump fifo_csv_dumper_1232;
    csv_file_dump cstatus_csv_dumper_1232;
    df_fifo_monitor fifo_monitor_1232;
    df_fifo_intf fifo_intf_1233(clock,reset);
    assign fifo_intf_1233.rd_en = AESL_inst_myproject.layer2_out_1232_U.if_read & AESL_inst_myproject.layer2_out_1232_U.if_empty_n;
    assign fifo_intf_1233.wr_en = AESL_inst_myproject.layer2_out_1232_U.if_write & AESL_inst_myproject.layer2_out_1232_U.if_full_n;
    assign fifo_intf_1233.fifo_rd_block = 0;
    assign fifo_intf_1233.fifo_wr_block = 0;
    assign fifo_intf_1233.finish = finish;
    csv_file_dump fifo_csv_dumper_1233;
    csv_file_dump cstatus_csv_dumper_1233;
    df_fifo_monitor fifo_monitor_1233;
    df_fifo_intf fifo_intf_1234(clock,reset);
    assign fifo_intf_1234.rd_en = AESL_inst_myproject.layer2_out_1233_U.if_read & AESL_inst_myproject.layer2_out_1233_U.if_empty_n;
    assign fifo_intf_1234.wr_en = AESL_inst_myproject.layer2_out_1233_U.if_write & AESL_inst_myproject.layer2_out_1233_U.if_full_n;
    assign fifo_intf_1234.fifo_rd_block = 0;
    assign fifo_intf_1234.fifo_wr_block = 0;
    assign fifo_intf_1234.finish = finish;
    csv_file_dump fifo_csv_dumper_1234;
    csv_file_dump cstatus_csv_dumper_1234;
    df_fifo_monitor fifo_monitor_1234;
    df_fifo_intf fifo_intf_1235(clock,reset);
    assign fifo_intf_1235.rd_en = AESL_inst_myproject.layer2_out_1234_U.if_read & AESL_inst_myproject.layer2_out_1234_U.if_empty_n;
    assign fifo_intf_1235.wr_en = AESL_inst_myproject.layer2_out_1234_U.if_write & AESL_inst_myproject.layer2_out_1234_U.if_full_n;
    assign fifo_intf_1235.fifo_rd_block = 0;
    assign fifo_intf_1235.fifo_wr_block = 0;
    assign fifo_intf_1235.finish = finish;
    csv_file_dump fifo_csv_dumper_1235;
    csv_file_dump cstatus_csv_dumper_1235;
    df_fifo_monitor fifo_monitor_1235;
    df_fifo_intf fifo_intf_1236(clock,reset);
    assign fifo_intf_1236.rd_en = AESL_inst_myproject.layer2_out_1235_U.if_read & AESL_inst_myproject.layer2_out_1235_U.if_empty_n;
    assign fifo_intf_1236.wr_en = AESL_inst_myproject.layer2_out_1235_U.if_write & AESL_inst_myproject.layer2_out_1235_U.if_full_n;
    assign fifo_intf_1236.fifo_rd_block = 0;
    assign fifo_intf_1236.fifo_wr_block = 0;
    assign fifo_intf_1236.finish = finish;
    csv_file_dump fifo_csv_dumper_1236;
    csv_file_dump cstatus_csv_dumper_1236;
    df_fifo_monitor fifo_monitor_1236;
    df_fifo_intf fifo_intf_1237(clock,reset);
    assign fifo_intf_1237.rd_en = AESL_inst_myproject.layer2_out_1236_U.if_read & AESL_inst_myproject.layer2_out_1236_U.if_empty_n;
    assign fifo_intf_1237.wr_en = AESL_inst_myproject.layer2_out_1236_U.if_write & AESL_inst_myproject.layer2_out_1236_U.if_full_n;
    assign fifo_intf_1237.fifo_rd_block = 0;
    assign fifo_intf_1237.fifo_wr_block = 0;
    assign fifo_intf_1237.finish = finish;
    csv_file_dump fifo_csv_dumper_1237;
    csv_file_dump cstatus_csv_dumper_1237;
    df_fifo_monitor fifo_monitor_1237;
    df_fifo_intf fifo_intf_1238(clock,reset);
    assign fifo_intf_1238.rd_en = AESL_inst_myproject.layer2_out_1237_U.if_read & AESL_inst_myproject.layer2_out_1237_U.if_empty_n;
    assign fifo_intf_1238.wr_en = AESL_inst_myproject.layer2_out_1237_U.if_write & AESL_inst_myproject.layer2_out_1237_U.if_full_n;
    assign fifo_intf_1238.fifo_rd_block = 0;
    assign fifo_intf_1238.fifo_wr_block = 0;
    assign fifo_intf_1238.finish = finish;
    csv_file_dump fifo_csv_dumper_1238;
    csv_file_dump cstatus_csv_dumper_1238;
    df_fifo_monitor fifo_monitor_1238;
    df_fifo_intf fifo_intf_1239(clock,reset);
    assign fifo_intf_1239.rd_en = AESL_inst_myproject.layer2_out_1238_U.if_read & AESL_inst_myproject.layer2_out_1238_U.if_empty_n;
    assign fifo_intf_1239.wr_en = AESL_inst_myproject.layer2_out_1238_U.if_write & AESL_inst_myproject.layer2_out_1238_U.if_full_n;
    assign fifo_intf_1239.fifo_rd_block = 0;
    assign fifo_intf_1239.fifo_wr_block = 0;
    assign fifo_intf_1239.finish = finish;
    csv_file_dump fifo_csv_dumper_1239;
    csv_file_dump cstatus_csv_dumper_1239;
    df_fifo_monitor fifo_monitor_1239;
    df_fifo_intf fifo_intf_1240(clock,reset);
    assign fifo_intf_1240.rd_en = AESL_inst_myproject.layer2_out_1239_U.if_read & AESL_inst_myproject.layer2_out_1239_U.if_empty_n;
    assign fifo_intf_1240.wr_en = AESL_inst_myproject.layer2_out_1239_U.if_write & AESL_inst_myproject.layer2_out_1239_U.if_full_n;
    assign fifo_intf_1240.fifo_rd_block = 0;
    assign fifo_intf_1240.fifo_wr_block = 0;
    assign fifo_intf_1240.finish = finish;
    csv_file_dump fifo_csv_dumper_1240;
    csv_file_dump cstatus_csv_dumper_1240;
    df_fifo_monitor fifo_monitor_1240;
    df_fifo_intf fifo_intf_1241(clock,reset);
    assign fifo_intf_1241.rd_en = AESL_inst_myproject.layer2_out_1240_U.if_read & AESL_inst_myproject.layer2_out_1240_U.if_empty_n;
    assign fifo_intf_1241.wr_en = AESL_inst_myproject.layer2_out_1240_U.if_write & AESL_inst_myproject.layer2_out_1240_U.if_full_n;
    assign fifo_intf_1241.fifo_rd_block = 0;
    assign fifo_intf_1241.fifo_wr_block = 0;
    assign fifo_intf_1241.finish = finish;
    csv_file_dump fifo_csv_dumper_1241;
    csv_file_dump cstatus_csv_dumper_1241;
    df_fifo_monitor fifo_monitor_1241;
    df_fifo_intf fifo_intf_1242(clock,reset);
    assign fifo_intf_1242.rd_en = AESL_inst_myproject.layer2_out_1241_U.if_read & AESL_inst_myproject.layer2_out_1241_U.if_empty_n;
    assign fifo_intf_1242.wr_en = AESL_inst_myproject.layer2_out_1241_U.if_write & AESL_inst_myproject.layer2_out_1241_U.if_full_n;
    assign fifo_intf_1242.fifo_rd_block = 0;
    assign fifo_intf_1242.fifo_wr_block = 0;
    assign fifo_intf_1242.finish = finish;
    csv_file_dump fifo_csv_dumper_1242;
    csv_file_dump cstatus_csv_dumper_1242;
    df_fifo_monitor fifo_monitor_1242;
    df_fifo_intf fifo_intf_1243(clock,reset);
    assign fifo_intf_1243.rd_en = AESL_inst_myproject.layer2_out_1242_U.if_read & AESL_inst_myproject.layer2_out_1242_U.if_empty_n;
    assign fifo_intf_1243.wr_en = AESL_inst_myproject.layer2_out_1242_U.if_write & AESL_inst_myproject.layer2_out_1242_U.if_full_n;
    assign fifo_intf_1243.fifo_rd_block = 0;
    assign fifo_intf_1243.fifo_wr_block = 0;
    assign fifo_intf_1243.finish = finish;
    csv_file_dump fifo_csv_dumper_1243;
    csv_file_dump cstatus_csv_dumper_1243;
    df_fifo_monitor fifo_monitor_1243;
    df_fifo_intf fifo_intf_1244(clock,reset);
    assign fifo_intf_1244.rd_en = AESL_inst_myproject.layer2_out_1243_U.if_read & AESL_inst_myproject.layer2_out_1243_U.if_empty_n;
    assign fifo_intf_1244.wr_en = AESL_inst_myproject.layer2_out_1243_U.if_write & AESL_inst_myproject.layer2_out_1243_U.if_full_n;
    assign fifo_intf_1244.fifo_rd_block = 0;
    assign fifo_intf_1244.fifo_wr_block = 0;
    assign fifo_intf_1244.finish = finish;
    csv_file_dump fifo_csv_dumper_1244;
    csv_file_dump cstatus_csv_dumper_1244;
    df_fifo_monitor fifo_monitor_1244;
    df_fifo_intf fifo_intf_1245(clock,reset);
    assign fifo_intf_1245.rd_en = AESL_inst_myproject.layer2_out_1244_U.if_read & AESL_inst_myproject.layer2_out_1244_U.if_empty_n;
    assign fifo_intf_1245.wr_en = AESL_inst_myproject.layer2_out_1244_U.if_write & AESL_inst_myproject.layer2_out_1244_U.if_full_n;
    assign fifo_intf_1245.fifo_rd_block = 0;
    assign fifo_intf_1245.fifo_wr_block = 0;
    assign fifo_intf_1245.finish = finish;
    csv_file_dump fifo_csv_dumper_1245;
    csv_file_dump cstatus_csv_dumper_1245;
    df_fifo_monitor fifo_monitor_1245;
    df_fifo_intf fifo_intf_1246(clock,reset);
    assign fifo_intf_1246.rd_en = AESL_inst_myproject.layer2_out_1245_U.if_read & AESL_inst_myproject.layer2_out_1245_U.if_empty_n;
    assign fifo_intf_1246.wr_en = AESL_inst_myproject.layer2_out_1245_U.if_write & AESL_inst_myproject.layer2_out_1245_U.if_full_n;
    assign fifo_intf_1246.fifo_rd_block = 0;
    assign fifo_intf_1246.fifo_wr_block = 0;
    assign fifo_intf_1246.finish = finish;
    csv_file_dump fifo_csv_dumper_1246;
    csv_file_dump cstatus_csv_dumper_1246;
    df_fifo_monitor fifo_monitor_1246;
    df_fifo_intf fifo_intf_1247(clock,reset);
    assign fifo_intf_1247.rd_en = AESL_inst_myproject.layer2_out_1246_U.if_read & AESL_inst_myproject.layer2_out_1246_U.if_empty_n;
    assign fifo_intf_1247.wr_en = AESL_inst_myproject.layer2_out_1246_U.if_write & AESL_inst_myproject.layer2_out_1246_U.if_full_n;
    assign fifo_intf_1247.fifo_rd_block = 0;
    assign fifo_intf_1247.fifo_wr_block = 0;
    assign fifo_intf_1247.finish = finish;
    csv_file_dump fifo_csv_dumper_1247;
    csv_file_dump cstatus_csv_dumper_1247;
    df_fifo_monitor fifo_monitor_1247;
    df_fifo_intf fifo_intf_1248(clock,reset);
    assign fifo_intf_1248.rd_en = AESL_inst_myproject.layer2_out_1247_U.if_read & AESL_inst_myproject.layer2_out_1247_U.if_empty_n;
    assign fifo_intf_1248.wr_en = AESL_inst_myproject.layer2_out_1247_U.if_write & AESL_inst_myproject.layer2_out_1247_U.if_full_n;
    assign fifo_intf_1248.fifo_rd_block = 0;
    assign fifo_intf_1248.fifo_wr_block = 0;
    assign fifo_intf_1248.finish = finish;
    csv_file_dump fifo_csv_dumper_1248;
    csv_file_dump cstatus_csv_dumper_1248;
    df_fifo_monitor fifo_monitor_1248;
    df_fifo_intf fifo_intf_1249(clock,reset);
    assign fifo_intf_1249.rd_en = AESL_inst_myproject.layer2_out_1248_U.if_read & AESL_inst_myproject.layer2_out_1248_U.if_empty_n;
    assign fifo_intf_1249.wr_en = AESL_inst_myproject.layer2_out_1248_U.if_write & AESL_inst_myproject.layer2_out_1248_U.if_full_n;
    assign fifo_intf_1249.fifo_rd_block = 0;
    assign fifo_intf_1249.fifo_wr_block = 0;
    assign fifo_intf_1249.finish = finish;
    csv_file_dump fifo_csv_dumper_1249;
    csv_file_dump cstatus_csv_dumper_1249;
    df_fifo_monitor fifo_monitor_1249;
    df_fifo_intf fifo_intf_1250(clock,reset);
    assign fifo_intf_1250.rd_en = AESL_inst_myproject.layer2_out_1249_U.if_read & AESL_inst_myproject.layer2_out_1249_U.if_empty_n;
    assign fifo_intf_1250.wr_en = AESL_inst_myproject.layer2_out_1249_U.if_write & AESL_inst_myproject.layer2_out_1249_U.if_full_n;
    assign fifo_intf_1250.fifo_rd_block = 0;
    assign fifo_intf_1250.fifo_wr_block = 0;
    assign fifo_intf_1250.finish = finish;
    csv_file_dump fifo_csv_dumper_1250;
    csv_file_dump cstatus_csv_dumper_1250;
    df_fifo_monitor fifo_monitor_1250;
    df_fifo_intf fifo_intf_1251(clock,reset);
    assign fifo_intf_1251.rd_en = AESL_inst_myproject.layer2_out_1250_U.if_read & AESL_inst_myproject.layer2_out_1250_U.if_empty_n;
    assign fifo_intf_1251.wr_en = AESL_inst_myproject.layer2_out_1250_U.if_write & AESL_inst_myproject.layer2_out_1250_U.if_full_n;
    assign fifo_intf_1251.fifo_rd_block = 0;
    assign fifo_intf_1251.fifo_wr_block = 0;
    assign fifo_intf_1251.finish = finish;
    csv_file_dump fifo_csv_dumper_1251;
    csv_file_dump cstatus_csv_dumper_1251;
    df_fifo_monitor fifo_monitor_1251;
    df_fifo_intf fifo_intf_1252(clock,reset);
    assign fifo_intf_1252.rd_en = AESL_inst_myproject.layer2_out_1251_U.if_read & AESL_inst_myproject.layer2_out_1251_U.if_empty_n;
    assign fifo_intf_1252.wr_en = AESL_inst_myproject.layer2_out_1251_U.if_write & AESL_inst_myproject.layer2_out_1251_U.if_full_n;
    assign fifo_intf_1252.fifo_rd_block = 0;
    assign fifo_intf_1252.fifo_wr_block = 0;
    assign fifo_intf_1252.finish = finish;
    csv_file_dump fifo_csv_dumper_1252;
    csv_file_dump cstatus_csv_dumper_1252;
    df_fifo_monitor fifo_monitor_1252;
    df_fifo_intf fifo_intf_1253(clock,reset);
    assign fifo_intf_1253.rd_en = AESL_inst_myproject.layer2_out_1252_U.if_read & AESL_inst_myproject.layer2_out_1252_U.if_empty_n;
    assign fifo_intf_1253.wr_en = AESL_inst_myproject.layer2_out_1252_U.if_write & AESL_inst_myproject.layer2_out_1252_U.if_full_n;
    assign fifo_intf_1253.fifo_rd_block = 0;
    assign fifo_intf_1253.fifo_wr_block = 0;
    assign fifo_intf_1253.finish = finish;
    csv_file_dump fifo_csv_dumper_1253;
    csv_file_dump cstatus_csv_dumper_1253;
    df_fifo_monitor fifo_monitor_1253;
    df_fifo_intf fifo_intf_1254(clock,reset);
    assign fifo_intf_1254.rd_en = AESL_inst_myproject.layer2_out_1253_U.if_read & AESL_inst_myproject.layer2_out_1253_U.if_empty_n;
    assign fifo_intf_1254.wr_en = AESL_inst_myproject.layer2_out_1253_U.if_write & AESL_inst_myproject.layer2_out_1253_U.if_full_n;
    assign fifo_intf_1254.fifo_rd_block = 0;
    assign fifo_intf_1254.fifo_wr_block = 0;
    assign fifo_intf_1254.finish = finish;
    csv_file_dump fifo_csv_dumper_1254;
    csv_file_dump cstatus_csv_dumper_1254;
    df_fifo_monitor fifo_monitor_1254;
    df_fifo_intf fifo_intf_1255(clock,reset);
    assign fifo_intf_1255.rd_en = AESL_inst_myproject.layer2_out_1254_U.if_read & AESL_inst_myproject.layer2_out_1254_U.if_empty_n;
    assign fifo_intf_1255.wr_en = AESL_inst_myproject.layer2_out_1254_U.if_write & AESL_inst_myproject.layer2_out_1254_U.if_full_n;
    assign fifo_intf_1255.fifo_rd_block = 0;
    assign fifo_intf_1255.fifo_wr_block = 0;
    assign fifo_intf_1255.finish = finish;
    csv_file_dump fifo_csv_dumper_1255;
    csv_file_dump cstatus_csv_dumper_1255;
    df_fifo_monitor fifo_monitor_1255;
    df_fifo_intf fifo_intf_1256(clock,reset);
    assign fifo_intf_1256.rd_en = AESL_inst_myproject.layer2_out_1255_U.if_read & AESL_inst_myproject.layer2_out_1255_U.if_empty_n;
    assign fifo_intf_1256.wr_en = AESL_inst_myproject.layer2_out_1255_U.if_write & AESL_inst_myproject.layer2_out_1255_U.if_full_n;
    assign fifo_intf_1256.fifo_rd_block = 0;
    assign fifo_intf_1256.fifo_wr_block = 0;
    assign fifo_intf_1256.finish = finish;
    csv_file_dump fifo_csv_dumper_1256;
    csv_file_dump cstatus_csv_dumper_1256;
    df_fifo_monitor fifo_monitor_1256;
    df_fifo_intf fifo_intf_1257(clock,reset);
    assign fifo_intf_1257.rd_en = AESL_inst_myproject.layer2_out_1256_U.if_read & AESL_inst_myproject.layer2_out_1256_U.if_empty_n;
    assign fifo_intf_1257.wr_en = AESL_inst_myproject.layer2_out_1256_U.if_write & AESL_inst_myproject.layer2_out_1256_U.if_full_n;
    assign fifo_intf_1257.fifo_rd_block = 0;
    assign fifo_intf_1257.fifo_wr_block = 0;
    assign fifo_intf_1257.finish = finish;
    csv_file_dump fifo_csv_dumper_1257;
    csv_file_dump cstatus_csv_dumper_1257;
    df_fifo_monitor fifo_monitor_1257;
    df_fifo_intf fifo_intf_1258(clock,reset);
    assign fifo_intf_1258.rd_en = AESL_inst_myproject.layer2_out_1257_U.if_read & AESL_inst_myproject.layer2_out_1257_U.if_empty_n;
    assign fifo_intf_1258.wr_en = AESL_inst_myproject.layer2_out_1257_U.if_write & AESL_inst_myproject.layer2_out_1257_U.if_full_n;
    assign fifo_intf_1258.fifo_rd_block = 0;
    assign fifo_intf_1258.fifo_wr_block = 0;
    assign fifo_intf_1258.finish = finish;
    csv_file_dump fifo_csv_dumper_1258;
    csv_file_dump cstatus_csv_dumper_1258;
    df_fifo_monitor fifo_monitor_1258;
    df_fifo_intf fifo_intf_1259(clock,reset);
    assign fifo_intf_1259.rd_en = AESL_inst_myproject.layer2_out_1258_U.if_read & AESL_inst_myproject.layer2_out_1258_U.if_empty_n;
    assign fifo_intf_1259.wr_en = AESL_inst_myproject.layer2_out_1258_U.if_write & AESL_inst_myproject.layer2_out_1258_U.if_full_n;
    assign fifo_intf_1259.fifo_rd_block = 0;
    assign fifo_intf_1259.fifo_wr_block = 0;
    assign fifo_intf_1259.finish = finish;
    csv_file_dump fifo_csv_dumper_1259;
    csv_file_dump cstatus_csv_dumper_1259;
    df_fifo_monitor fifo_monitor_1259;
    df_fifo_intf fifo_intf_1260(clock,reset);
    assign fifo_intf_1260.rd_en = AESL_inst_myproject.layer2_out_1259_U.if_read & AESL_inst_myproject.layer2_out_1259_U.if_empty_n;
    assign fifo_intf_1260.wr_en = AESL_inst_myproject.layer2_out_1259_U.if_write & AESL_inst_myproject.layer2_out_1259_U.if_full_n;
    assign fifo_intf_1260.fifo_rd_block = 0;
    assign fifo_intf_1260.fifo_wr_block = 0;
    assign fifo_intf_1260.finish = finish;
    csv_file_dump fifo_csv_dumper_1260;
    csv_file_dump cstatus_csv_dumper_1260;
    df_fifo_monitor fifo_monitor_1260;
    df_fifo_intf fifo_intf_1261(clock,reset);
    assign fifo_intf_1261.rd_en = AESL_inst_myproject.layer2_out_1260_U.if_read & AESL_inst_myproject.layer2_out_1260_U.if_empty_n;
    assign fifo_intf_1261.wr_en = AESL_inst_myproject.layer2_out_1260_U.if_write & AESL_inst_myproject.layer2_out_1260_U.if_full_n;
    assign fifo_intf_1261.fifo_rd_block = 0;
    assign fifo_intf_1261.fifo_wr_block = 0;
    assign fifo_intf_1261.finish = finish;
    csv_file_dump fifo_csv_dumper_1261;
    csv_file_dump cstatus_csv_dumper_1261;
    df_fifo_monitor fifo_monitor_1261;
    df_fifo_intf fifo_intf_1262(clock,reset);
    assign fifo_intf_1262.rd_en = AESL_inst_myproject.layer2_out_1261_U.if_read & AESL_inst_myproject.layer2_out_1261_U.if_empty_n;
    assign fifo_intf_1262.wr_en = AESL_inst_myproject.layer2_out_1261_U.if_write & AESL_inst_myproject.layer2_out_1261_U.if_full_n;
    assign fifo_intf_1262.fifo_rd_block = 0;
    assign fifo_intf_1262.fifo_wr_block = 0;
    assign fifo_intf_1262.finish = finish;
    csv_file_dump fifo_csv_dumper_1262;
    csv_file_dump cstatus_csv_dumper_1262;
    df_fifo_monitor fifo_monitor_1262;
    df_fifo_intf fifo_intf_1263(clock,reset);
    assign fifo_intf_1263.rd_en = AESL_inst_myproject.layer2_out_1262_U.if_read & AESL_inst_myproject.layer2_out_1262_U.if_empty_n;
    assign fifo_intf_1263.wr_en = AESL_inst_myproject.layer2_out_1262_U.if_write & AESL_inst_myproject.layer2_out_1262_U.if_full_n;
    assign fifo_intf_1263.fifo_rd_block = 0;
    assign fifo_intf_1263.fifo_wr_block = 0;
    assign fifo_intf_1263.finish = finish;
    csv_file_dump fifo_csv_dumper_1263;
    csv_file_dump cstatus_csv_dumper_1263;
    df_fifo_monitor fifo_monitor_1263;
    df_fifo_intf fifo_intf_1264(clock,reset);
    assign fifo_intf_1264.rd_en = AESL_inst_myproject.layer2_out_1263_U.if_read & AESL_inst_myproject.layer2_out_1263_U.if_empty_n;
    assign fifo_intf_1264.wr_en = AESL_inst_myproject.layer2_out_1263_U.if_write & AESL_inst_myproject.layer2_out_1263_U.if_full_n;
    assign fifo_intf_1264.fifo_rd_block = 0;
    assign fifo_intf_1264.fifo_wr_block = 0;
    assign fifo_intf_1264.finish = finish;
    csv_file_dump fifo_csv_dumper_1264;
    csv_file_dump cstatus_csv_dumper_1264;
    df_fifo_monitor fifo_monitor_1264;
    df_fifo_intf fifo_intf_1265(clock,reset);
    assign fifo_intf_1265.rd_en = AESL_inst_myproject.layer2_out_1264_U.if_read & AESL_inst_myproject.layer2_out_1264_U.if_empty_n;
    assign fifo_intf_1265.wr_en = AESL_inst_myproject.layer2_out_1264_U.if_write & AESL_inst_myproject.layer2_out_1264_U.if_full_n;
    assign fifo_intf_1265.fifo_rd_block = 0;
    assign fifo_intf_1265.fifo_wr_block = 0;
    assign fifo_intf_1265.finish = finish;
    csv_file_dump fifo_csv_dumper_1265;
    csv_file_dump cstatus_csv_dumper_1265;
    df_fifo_monitor fifo_monitor_1265;
    df_fifo_intf fifo_intf_1266(clock,reset);
    assign fifo_intf_1266.rd_en = AESL_inst_myproject.layer2_out_1265_U.if_read & AESL_inst_myproject.layer2_out_1265_U.if_empty_n;
    assign fifo_intf_1266.wr_en = AESL_inst_myproject.layer2_out_1265_U.if_write & AESL_inst_myproject.layer2_out_1265_U.if_full_n;
    assign fifo_intf_1266.fifo_rd_block = 0;
    assign fifo_intf_1266.fifo_wr_block = 0;
    assign fifo_intf_1266.finish = finish;
    csv_file_dump fifo_csv_dumper_1266;
    csv_file_dump cstatus_csv_dumper_1266;
    df_fifo_monitor fifo_monitor_1266;
    df_fifo_intf fifo_intf_1267(clock,reset);
    assign fifo_intf_1267.rd_en = AESL_inst_myproject.layer2_out_1266_U.if_read & AESL_inst_myproject.layer2_out_1266_U.if_empty_n;
    assign fifo_intf_1267.wr_en = AESL_inst_myproject.layer2_out_1266_U.if_write & AESL_inst_myproject.layer2_out_1266_U.if_full_n;
    assign fifo_intf_1267.fifo_rd_block = 0;
    assign fifo_intf_1267.fifo_wr_block = 0;
    assign fifo_intf_1267.finish = finish;
    csv_file_dump fifo_csv_dumper_1267;
    csv_file_dump cstatus_csv_dumper_1267;
    df_fifo_monitor fifo_monitor_1267;
    df_fifo_intf fifo_intf_1268(clock,reset);
    assign fifo_intf_1268.rd_en = AESL_inst_myproject.layer2_out_1267_U.if_read & AESL_inst_myproject.layer2_out_1267_U.if_empty_n;
    assign fifo_intf_1268.wr_en = AESL_inst_myproject.layer2_out_1267_U.if_write & AESL_inst_myproject.layer2_out_1267_U.if_full_n;
    assign fifo_intf_1268.fifo_rd_block = 0;
    assign fifo_intf_1268.fifo_wr_block = 0;
    assign fifo_intf_1268.finish = finish;
    csv_file_dump fifo_csv_dumper_1268;
    csv_file_dump cstatus_csv_dumper_1268;
    df_fifo_monitor fifo_monitor_1268;
    df_fifo_intf fifo_intf_1269(clock,reset);
    assign fifo_intf_1269.rd_en = AESL_inst_myproject.layer2_out_1268_U.if_read & AESL_inst_myproject.layer2_out_1268_U.if_empty_n;
    assign fifo_intf_1269.wr_en = AESL_inst_myproject.layer2_out_1268_U.if_write & AESL_inst_myproject.layer2_out_1268_U.if_full_n;
    assign fifo_intf_1269.fifo_rd_block = 0;
    assign fifo_intf_1269.fifo_wr_block = 0;
    assign fifo_intf_1269.finish = finish;
    csv_file_dump fifo_csv_dumper_1269;
    csv_file_dump cstatus_csv_dumper_1269;
    df_fifo_monitor fifo_monitor_1269;
    df_fifo_intf fifo_intf_1270(clock,reset);
    assign fifo_intf_1270.rd_en = AESL_inst_myproject.layer2_out_1269_U.if_read & AESL_inst_myproject.layer2_out_1269_U.if_empty_n;
    assign fifo_intf_1270.wr_en = AESL_inst_myproject.layer2_out_1269_U.if_write & AESL_inst_myproject.layer2_out_1269_U.if_full_n;
    assign fifo_intf_1270.fifo_rd_block = 0;
    assign fifo_intf_1270.fifo_wr_block = 0;
    assign fifo_intf_1270.finish = finish;
    csv_file_dump fifo_csv_dumper_1270;
    csv_file_dump cstatus_csv_dumper_1270;
    df_fifo_monitor fifo_monitor_1270;
    df_fifo_intf fifo_intf_1271(clock,reset);
    assign fifo_intf_1271.rd_en = AESL_inst_myproject.layer2_out_1270_U.if_read & AESL_inst_myproject.layer2_out_1270_U.if_empty_n;
    assign fifo_intf_1271.wr_en = AESL_inst_myproject.layer2_out_1270_U.if_write & AESL_inst_myproject.layer2_out_1270_U.if_full_n;
    assign fifo_intf_1271.fifo_rd_block = 0;
    assign fifo_intf_1271.fifo_wr_block = 0;
    assign fifo_intf_1271.finish = finish;
    csv_file_dump fifo_csv_dumper_1271;
    csv_file_dump cstatus_csv_dumper_1271;
    df_fifo_monitor fifo_monitor_1271;
    df_fifo_intf fifo_intf_1272(clock,reset);
    assign fifo_intf_1272.rd_en = AESL_inst_myproject.layer2_out_1271_U.if_read & AESL_inst_myproject.layer2_out_1271_U.if_empty_n;
    assign fifo_intf_1272.wr_en = AESL_inst_myproject.layer2_out_1271_U.if_write & AESL_inst_myproject.layer2_out_1271_U.if_full_n;
    assign fifo_intf_1272.fifo_rd_block = 0;
    assign fifo_intf_1272.fifo_wr_block = 0;
    assign fifo_intf_1272.finish = finish;
    csv_file_dump fifo_csv_dumper_1272;
    csv_file_dump cstatus_csv_dumper_1272;
    df_fifo_monitor fifo_monitor_1272;
    df_fifo_intf fifo_intf_1273(clock,reset);
    assign fifo_intf_1273.rd_en = AESL_inst_myproject.layer2_out_1272_U.if_read & AESL_inst_myproject.layer2_out_1272_U.if_empty_n;
    assign fifo_intf_1273.wr_en = AESL_inst_myproject.layer2_out_1272_U.if_write & AESL_inst_myproject.layer2_out_1272_U.if_full_n;
    assign fifo_intf_1273.fifo_rd_block = 0;
    assign fifo_intf_1273.fifo_wr_block = 0;
    assign fifo_intf_1273.finish = finish;
    csv_file_dump fifo_csv_dumper_1273;
    csv_file_dump cstatus_csv_dumper_1273;
    df_fifo_monitor fifo_monitor_1273;
    df_fifo_intf fifo_intf_1274(clock,reset);
    assign fifo_intf_1274.rd_en = AESL_inst_myproject.layer2_out_1273_U.if_read & AESL_inst_myproject.layer2_out_1273_U.if_empty_n;
    assign fifo_intf_1274.wr_en = AESL_inst_myproject.layer2_out_1273_U.if_write & AESL_inst_myproject.layer2_out_1273_U.if_full_n;
    assign fifo_intf_1274.fifo_rd_block = 0;
    assign fifo_intf_1274.fifo_wr_block = 0;
    assign fifo_intf_1274.finish = finish;
    csv_file_dump fifo_csv_dumper_1274;
    csv_file_dump cstatus_csv_dumper_1274;
    df_fifo_monitor fifo_monitor_1274;
    df_fifo_intf fifo_intf_1275(clock,reset);
    assign fifo_intf_1275.rd_en = AESL_inst_myproject.layer2_out_1274_U.if_read & AESL_inst_myproject.layer2_out_1274_U.if_empty_n;
    assign fifo_intf_1275.wr_en = AESL_inst_myproject.layer2_out_1274_U.if_write & AESL_inst_myproject.layer2_out_1274_U.if_full_n;
    assign fifo_intf_1275.fifo_rd_block = 0;
    assign fifo_intf_1275.fifo_wr_block = 0;
    assign fifo_intf_1275.finish = finish;
    csv_file_dump fifo_csv_dumper_1275;
    csv_file_dump cstatus_csv_dumper_1275;
    df_fifo_monitor fifo_monitor_1275;
    df_fifo_intf fifo_intf_1276(clock,reset);
    assign fifo_intf_1276.rd_en = AESL_inst_myproject.layer2_out_1275_U.if_read & AESL_inst_myproject.layer2_out_1275_U.if_empty_n;
    assign fifo_intf_1276.wr_en = AESL_inst_myproject.layer2_out_1275_U.if_write & AESL_inst_myproject.layer2_out_1275_U.if_full_n;
    assign fifo_intf_1276.fifo_rd_block = 0;
    assign fifo_intf_1276.fifo_wr_block = 0;
    assign fifo_intf_1276.finish = finish;
    csv_file_dump fifo_csv_dumper_1276;
    csv_file_dump cstatus_csv_dumper_1276;
    df_fifo_monitor fifo_monitor_1276;
    df_fifo_intf fifo_intf_1277(clock,reset);
    assign fifo_intf_1277.rd_en = AESL_inst_myproject.layer2_out_1276_U.if_read & AESL_inst_myproject.layer2_out_1276_U.if_empty_n;
    assign fifo_intf_1277.wr_en = AESL_inst_myproject.layer2_out_1276_U.if_write & AESL_inst_myproject.layer2_out_1276_U.if_full_n;
    assign fifo_intf_1277.fifo_rd_block = 0;
    assign fifo_intf_1277.fifo_wr_block = 0;
    assign fifo_intf_1277.finish = finish;
    csv_file_dump fifo_csv_dumper_1277;
    csv_file_dump cstatus_csv_dumper_1277;
    df_fifo_monitor fifo_monitor_1277;
    df_fifo_intf fifo_intf_1278(clock,reset);
    assign fifo_intf_1278.rd_en = AESL_inst_myproject.layer2_out_1277_U.if_read & AESL_inst_myproject.layer2_out_1277_U.if_empty_n;
    assign fifo_intf_1278.wr_en = AESL_inst_myproject.layer2_out_1277_U.if_write & AESL_inst_myproject.layer2_out_1277_U.if_full_n;
    assign fifo_intf_1278.fifo_rd_block = 0;
    assign fifo_intf_1278.fifo_wr_block = 0;
    assign fifo_intf_1278.finish = finish;
    csv_file_dump fifo_csv_dumper_1278;
    csv_file_dump cstatus_csv_dumper_1278;
    df_fifo_monitor fifo_monitor_1278;
    df_fifo_intf fifo_intf_1279(clock,reset);
    assign fifo_intf_1279.rd_en = AESL_inst_myproject.layer2_out_1278_U.if_read & AESL_inst_myproject.layer2_out_1278_U.if_empty_n;
    assign fifo_intf_1279.wr_en = AESL_inst_myproject.layer2_out_1278_U.if_write & AESL_inst_myproject.layer2_out_1278_U.if_full_n;
    assign fifo_intf_1279.fifo_rd_block = 0;
    assign fifo_intf_1279.fifo_wr_block = 0;
    assign fifo_intf_1279.finish = finish;
    csv_file_dump fifo_csv_dumper_1279;
    csv_file_dump cstatus_csv_dumper_1279;
    df_fifo_monitor fifo_monitor_1279;
    df_fifo_intf fifo_intf_1280(clock,reset);
    assign fifo_intf_1280.rd_en = AESL_inst_myproject.layer2_out_1279_U.if_read & AESL_inst_myproject.layer2_out_1279_U.if_empty_n;
    assign fifo_intf_1280.wr_en = AESL_inst_myproject.layer2_out_1279_U.if_write & AESL_inst_myproject.layer2_out_1279_U.if_full_n;
    assign fifo_intf_1280.fifo_rd_block = 0;
    assign fifo_intf_1280.fifo_wr_block = 0;
    assign fifo_intf_1280.finish = finish;
    csv_file_dump fifo_csv_dumper_1280;
    csv_file_dump cstatus_csv_dumper_1280;
    df_fifo_monitor fifo_monitor_1280;
    df_fifo_intf fifo_intf_1281(clock,reset);
    assign fifo_intf_1281.rd_en = AESL_inst_myproject.layer2_out_1280_U.if_read & AESL_inst_myproject.layer2_out_1280_U.if_empty_n;
    assign fifo_intf_1281.wr_en = AESL_inst_myproject.layer2_out_1280_U.if_write & AESL_inst_myproject.layer2_out_1280_U.if_full_n;
    assign fifo_intf_1281.fifo_rd_block = 0;
    assign fifo_intf_1281.fifo_wr_block = 0;
    assign fifo_intf_1281.finish = finish;
    csv_file_dump fifo_csv_dumper_1281;
    csv_file_dump cstatus_csv_dumper_1281;
    df_fifo_monitor fifo_monitor_1281;
    df_fifo_intf fifo_intf_1282(clock,reset);
    assign fifo_intf_1282.rd_en = AESL_inst_myproject.layer2_out_1281_U.if_read & AESL_inst_myproject.layer2_out_1281_U.if_empty_n;
    assign fifo_intf_1282.wr_en = AESL_inst_myproject.layer2_out_1281_U.if_write & AESL_inst_myproject.layer2_out_1281_U.if_full_n;
    assign fifo_intf_1282.fifo_rd_block = 0;
    assign fifo_intf_1282.fifo_wr_block = 0;
    assign fifo_intf_1282.finish = finish;
    csv_file_dump fifo_csv_dumper_1282;
    csv_file_dump cstatus_csv_dumper_1282;
    df_fifo_monitor fifo_monitor_1282;
    df_fifo_intf fifo_intf_1283(clock,reset);
    assign fifo_intf_1283.rd_en = AESL_inst_myproject.layer2_out_1282_U.if_read & AESL_inst_myproject.layer2_out_1282_U.if_empty_n;
    assign fifo_intf_1283.wr_en = AESL_inst_myproject.layer2_out_1282_U.if_write & AESL_inst_myproject.layer2_out_1282_U.if_full_n;
    assign fifo_intf_1283.fifo_rd_block = 0;
    assign fifo_intf_1283.fifo_wr_block = 0;
    assign fifo_intf_1283.finish = finish;
    csv_file_dump fifo_csv_dumper_1283;
    csv_file_dump cstatus_csv_dumper_1283;
    df_fifo_monitor fifo_monitor_1283;
    df_fifo_intf fifo_intf_1284(clock,reset);
    assign fifo_intf_1284.rd_en = AESL_inst_myproject.layer2_out_1283_U.if_read & AESL_inst_myproject.layer2_out_1283_U.if_empty_n;
    assign fifo_intf_1284.wr_en = AESL_inst_myproject.layer2_out_1283_U.if_write & AESL_inst_myproject.layer2_out_1283_U.if_full_n;
    assign fifo_intf_1284.fifo_rd_block = 0;
    assign fifo_intf_1284.fifo_wr_block = 0;
    assign fifo_intf_1284.finish = finish;
    csv_file_dump fifo_csv_dumper_1284;
    csv_file_dump cstatus_csv_dumper_1284;
    df_fifo_monitor fifo_monitor_1284;
    df_fifo_intf fifo_intf_1285(clock,reset);
    assign fifo_intf_1285.rd_en = AESL_inst_myproject.layer2_out_1284_U.if_read & AESL_inst_myproject.layer2_out_1284_U.if_empty_n;
    assign fifo_intf_1285.wr_en = AESL_inst_myproject.layer2_out_1284_U.if_write & AESL_inst_myproject.layer2_out_1284_U.if_full_n;
    assign fifo_intf_1285.fifo_rd_block = 0;
    assign fifo_intf_1285.fifo_wr_block = 0;
    assign fifo_intf_1285.finish = finish;
    csv_file_dump fifo_csv_dumper_1285;
    csv_file_dump cstatus_csv_dumper_1285;
    df_fifo_monitor fifo_monitor_1285;
    df_fifo_intf fifo_intf_1286(clock,reset);
    assign fifo_intf_1286.rd_en = AESL_inst_myproject.layer2_out_1285_U.if_read & AESL_inst_myproject.layer2_out_1285_U.if_empty_n;
    assign fifo_intf_1286.wr_en = AESL_inst_myproject.layer2_out_1285_U.if_write & AESL_inst_myproject.layer2_out_1285_U.if_full_n;
    assign fifo_intf_1286.fifo_rd_block = 0;
    assign fifo_intf_1286.fifo_wr_block = 0;
    assign fifo_intf_1286.finish = finish;
    csv_file_dump fifo_csv_dumper_1286;
    csv_file_dump cstatus_csv_dumper_1286;
    df_fifo_monitor fifo_monitor_1286;
    df_fifo_intf fifo_intf_1287(clock,reset);
    assign fifo_intf_1287.rd_en = AESL_inst_myproject.layer2_out_1286_U.if_read & AESL_inst_myproject.layer2_out_1286_U.if_empty_n;
    assign fifo_intf_1287.wr_en = AESL_inst_myproject.layer2_out_1286_U.if_write & AESL_inst_myproject.layer2_out_1286_U.if_full_n;
    assign fifo_intf_1287.fifo_rd_block = 0;
    assign fifo_intf_1287.fifo_wr_block = 0;
    assign fifo_intf_1287.finish = finish;
    csv_file_dump fifo_csv_dumper_1287;
    csv_file_dump cstatus_csv_dumper_1287;
    df_fifo_monitor fifo_monitor_1287;
    df_fifo_intf fifo_intf_1288(clock,reset);
    assign fifo_intf_1288.rd_en = AESL_inst_myproject.layer2_out_1287_U.if_read & AESL_inst_myproject.layer2_out_1287_U.if_empty_n;
    assign fifo_intf_1288.wr_en = AESL_inst_myproject.layer2_out_1287_U.if_write & AESL_inst_myproject.layer2_out_1287_U.if_full_n;
    assign fifo_intf_1288.fifo_rd_block = 0;
    assign fifo_intf_1288.fifo_wr_block = 0;
    assign fifo_intf_1288.finish = finish;
    csv_file_dump fifo_csv_dumper_1288;
    csv_file_dump cstatus_csv_dumper_1288;
    df_fifo_monitor fifo_monitor_1288;
    df_fifo_intf fifo_intf_1289(clock,reset);
    assign fifo_intf_1289.rd_en = AESL_inst_myproject.layer2_out_1288_U.if_read & AESL_inst_myproject.layer2_out_1288_U.if_empty_n;
    assign fifo_intf_1289.wr_en = AESL_inst_myproject.layer2_out_1288_U.if_write & AESL_inst_myproject.layer2_out_1288_U.if_full_n;
    assign fifo_intf_1289.fifo_rd_block = 0;
    assign fifo_intf_1289.fifo_wr_block = 0;
    assign fifo_intf_1289.finish = finish;
    csv_file_dump fifo_csv_dumper_1289;
    csv_file_dump cstatus_csv_dumper_1289;
    df_fifo_monitor fifo_monitor_1289;
    df_fifo_intf fifo_intf_1290(clock,reset);
    assign fifo_intf_1290.rd_en = AESL_inst_myproject.layer2_out_1289_U.if_read & AESL_inst_myproject.layer2_out_1289_U.if_empty_n;
    assign fifo_intf_1290.wr_en = AESL_inst_myproject.layer2_out_1289_U.if_write & AESL_inst_myproject.layer2_out_1289_U.if_full_n;
    assign fifo_intf_1290.fifo_rd_block = 0;
    assign fifo_intf_1290.fifo_wr_block = 0;
    assign fifo_intf_1290.finish = finish;
    csv_file_dump fifo_csv_dumper_1290;
    csv_file_dump cstatus_csv_dumper_1290;
    df_fifo_monitor fifo_monitor_1290;
    df_fifo_intf fifo_intf_1291(clock,reset);
    assign fifo_intf_1291.rd_en = AESL_inst_myproject.layer2_out_1290_U.if_read & AESL_inst_myproject.layer2_out_1290_U.if_empty_n;
    assign fifo_intf_1291.wr_en = AESL_inst_myproject.layer2_out_1290_U.if_write & AESL_inst_myproject.layer2_out_1290_U.if_full_n;
    assign fifo_intf_1291.fifo_rd_block = 0;
    assign fifo_intf_1291.fifo_wr_block = 0;
    assign fifo_intf_1291.finish = finish;
    csv_file_dump fifo_csv_dumper_1291;
    csv_file_dump cstatus_csv_dumper_1291;
    df_fifo_monitor fifo_monitor_1291;
    df_fifo_intf fifo_intf_1292(clock,reset);
    assign fifo_intf_1292.rd_en = AESL_inst_myproject.layer2_out_1291_U.if_read & AESL_inst_myproject.layer2_out_1291_U.if_empty_n;
    assign fifo_intf_1292.wr_en = AESL_inst_myproject.layer2_out_1291_U.if_write & AESL_inst_myproject.layer2_out_1291_U.if_full_n;
    assign fifo_intf_1292.fifo_rd_block = 0;
    assign fifo_intf_1292.fifo_wr_block = 0;
    assign fifo_intf_1292.finish = finish;
    csv_file_dump fifo_csv_dumper_1292;
    csv_file_dump cstatus_csv_dumper_1292;
    df_fifo_monitor fifo_monitor_1292;
    df_fifo_intf fifo_intf_1293(clock,reset);
    assign fifo_intf_1293.rd_en = AESL_inst_myproject.layer2_out_1292_U.if_read & AESL_inst_myproject.layer2_out_1292_U.if_empty_n;
    assign fifo_intf_1293.wr_en = AESL_inst_myproject.layer2_out_1292_U.if_write & AESL_inst_myproject.layer2_out_1292_U.if_full_n;
    assign fifo_intf_1293.fifo_rd_block = 0;
    assign fifo_intf_1293.fifo_wr_block = 0;
    assign fifo_intf_1293.finish = finish;
    csv_file_dump fifo_csv_dumper_1293;
    csv_file_dump cstatus_csv_dumper_1293;
    df_fifo_monitor fifo_monitor_1293;
    df_fifo_intf fifo_intf_1294(clock,reset);
    assign fifo_intf_1294.rd_en = AESL_inst_myproject.layer2_out_1293_U.if_read & AESL_inst_myproject.layer2_out_1293_U.if_empty_n;
    assign fifo_intf_1294.wr_en = AESL_inst_myproject.layer2_out_1293_U.if_write & AESL_inst_myproject.layer2_out_1293_U.if_full_n;
    assign fifo_intf_1294.fifo_rd_block = 0;
    assign fifo_intf_1294.fifo_wr_block = 0;
    assign fifo_intf_1294.finish = finish;
    csv_file_dump fifo_csv_dumper_1294;
    csv_file_dump cstatus_csv_dumper_1294;
    df_fifo_monitor fifo_monitor_1294;
    df_fifo_intf fifo_intf_1295(clock,reset);
    assign fifo_intf_1295.rd_en = AESL_inst_myproject.layer2_out_1294_U.if_read & AESL_inst_myproject.layer2_out_1294_U.if_empty_n;
    assign fifo_intf_1295.wr_en = AESL_inst_myproject.layer2_out_1294_U.if_write & AESL_inst_myproject.layer2_out_1294_U.if_full_n;
    assign fifo_intf_1295.fifo_rd_block = 0;
    assign fifo_intf_1295.fifo_wr_block = 0;
    assign fifo_intf_1295.finish = finish;
    csv_file_dump fifo_csv_dumper_1295;
    csv_file_dump cstatus_csv_dumper_1295;
    df_fifo_monitor fifo_monitor_1295;
    df_fifo_intf fifo_intf_1296(clock,reset);
    assign fifo_intf_1296.rd_en = AESL_inst_myproject.layer2_out_1295_U.if_read & AESL_inst_myproject.layer2_out_1295_U.if_empty_n;
    assign fifo_intf_1296.wr_en = AESL_inst_myproject.layer2_out_1295_U.if_write & AESL_inst_myproject.layer2_out_1295_U.if_full_n;
    assign fifo_intf_1296.fifo_rd_block = 0;
    assign fifo_intf_1296.fifo_wr_block = 0;
    assign fifo_intf_1296.finish = finish;
    csv_file_dump fifo_csv_dumper_1296;
    csv_file_dump cstatus_csv_dumper_1296;
    df_fifo_monitor fifo_monitor_1296;
    df_fifo_intf fifo_intf_1297(clock,reset);
    assign fifo_intf_1297.rd_en = AESL_inst_myproject.layer2_out_1296_U.if_read & AESL_inst_myproject.layer2_out_1296_U.if_empty_n;
    assign fifo_intf_1297.wr_en = AESL_inst_myproject.layer2_out_1296_U.if_write & AESL_inst_myproject.layer2_out_1296_U.if_full_n;
    assign fifo_intf_1297.fifo_rd_block = 0;
    assign fifo_intf_1297.fifo_wr_block = 0;
    assign fifo_intf_1297.finish = finish;
    csv_file_dump fifo_csv_dumper_1297;
    csv_file_dump cstatus_csv_dumper_1297;
    df_fifo_monitor fifo_monitor_1297;
    df_fifo_intf fifo_intf_1298(clock,reset);
    assign fifo_intf_1298.rd_en = AESL_inst_myproject.layer2_out_1297_U.if_read & AESL_inst_myproject.layer2_out_1297_U.if_empty_n;
    assign fifo_intf_1298.wr_en = AESL_inst_myproject.layer2_out_1297_U.if_write & AESL_inst_myproject.layer2_out_1297_U.if_full_n;
    assign fifo_intf_1298.fifo_rd_block = 0;
    assign fifo_intf_1298.fifo_wr_block = 0;
    assign fifo_intf_1298.finish = finish;
    csv_file_dump fifo_csv_dumper_1298;
    csv_file_dump cstatus_csv_dumper_1298;
    df_fifo_monitor fifo_monitor_1298;
    df_fifo_intf fifo_intf_1299(clock,reset);
    assign fifo_intf_1299.rd_en = AESL_inst_myproject.layer2_out_1298_U.if_read & AESL_inst_myproject.layer2_out_1298_U.if_empty_n;
    assign fifo_intf_1299.wr_en = AESL_inst_myproject.layer2_out_1298_U.if_write & AESL_inst_myproject.layer2_out_1298_U.if_full_n;
    assign fifo_intf_1299.fifo_rd_block = 0;
    assign fifo_intf_1299.fifo_wr_block = 0;
    assign fifo_intf_1299.finish = finish;
    csv_file_dump fifo_csv_dumper_1299;
    csv_file_dump cstatus_csv_dumper_1299;
    df_fifo_monitor fifo_monitor_1299;
    df_fifo_intf fifo_intf_1300(clock,reset);
    assign fifo_intf_1300.rd_en = AESL_inst_myproject.layer2_out_1299_U.if_read & AESL_inst_myproject.layer2_out_1299_U.if_empty_n;
    assign fifo_intf_1300.wr_en = AESL_inst_myproject.layer2_out_1299_U.if_write & AESL_inst_myproject.layer2_out_1299_U.if_full_n;
    assign fifo_intf_1300.fifo_rd_block = 0;
    assign fifo_intf_1300.fifo_wr_block = 0;
    assign fifo_intf_1300.finish = finish;
    csv_file_dump fifo_csv_dumper_1300;
    csv_file_dump cstatus_csv_dumper_1300;
    df_fifo_monitor fifo_monitor_1300;
    df_fifo_intf fifo_intf_1301(clock,reset);
    assign fifo_intf_1301.rd_en = AESL_inst_myproject.layer2_out_1300_U.if_read & AESL_inst_myproject.layer2_out_1300_U.if_empty_n;
    assign fifo_intf_1301.wr_en = AESL_inst_myproject.layer2_out_1300_U.if_write & AESL_inst_myproject.layer2_out_1300_U.if_full_n;
    assign fifo_intf_1301.fifo_rd_block = 0;
    assign fifo_intf_1301.fifo_wr_block = 0;
    assign fifo_intf_1301.finish = finish;
    csv_file_dump fifo_csv_dumper_1301;
    csv_file_dump cstatus_csv_dumper_1301;
    df_fifo_monitor fifo_monitor_1301;
    df_fifo_intf fifo_intf_1302(clock,reset);
    assign fifo_intf_1302.rd_en = AESL_inst_myproject.layer2_out_1301_U.if_read & AESL_inst_myproject.layer2_out_1301_U.if_empty_n;
    assign fifo_intf_1302.wr_en = AESL_inst_myproject.layer2_out_1301_U.if_write & AESL_inst_myproject.layer2_out_1301_U.if_full_n;
    assign fifo_intf_1302.fifo_rd_block = 0;
    assign fifo_intf_1302.fifo_wr_block = 0;
    assign fifo_intf_1302.finish = finish;
    csv_file_dump fifo_csv_dumper_1302;
    csv_file_dump cstatus_csv_dumper_1302;
    df_fifo_monitor fifo_monitor_1302;
    df_fifo_intf fifo_intf_1303(clock,reset);
    assign fifo_intf_1303.rd_en = AESL_inst_myproject.layer2_out_1302_U.if_read & AESL_inst_myproject.layer2_out_1302_U.if_empty_n;
    assign fifo_intf_1303.wr_en = AESL_inst_myproject.layer2_out_1302_U.if_write & AESL_inst_myproject.layer2_out_1302_U.if_full_n;
    assign fifo_intf_1303.fifo_rd_block = 0;
    assign fifo_intf_1303.fifo_wr_block = 0;
    assign fifo_intf_1303.finish = finish;
    csv_file_dump fifo_csv_dumper_1303;
    csv_file_dump cstatus_csv_dumper_1303;
    df_fifo_monitor fifo_monitor_1303;
    df_fifo_intf fifo_intf_1304(clock,reset);
    assign fifo_intf_1304.rd_en = AESL_inst_myproject.layer2_out_1303_U.if_read & AESL_inst_myproject.layer2_out_1303_U.if_empty_n;
    assign fifo_intf_1304.wr_en = AESL_inst_myproject.layer2_out_1303_U.if_write & AESL_inst_myproject.layer2_out_1303_U.if_full_n;
    assign fifo_intf_1304.fifo_rd_block = 0;
    assign fifo_intf_1304.fifo_wr_block = 0;
    assign fifo_intf_1304.finish = finish;
    csv_file_dump fifo_csv_dumper_1304;
    csv_file_dump cstatus_csv_dumper_1304;
    df_fifo_monitor fifo_monitor_1304;
    df_fifo_intf fifo_intf_1305(clock,reset);
    assign fifo_intf_1305.rd_en = AESL_inst_myproject.layer2_out_1304_U.if_read & AESL_inst_myproject.layer2_out_1304_U.if_empty_n;
    assign fifo_intf_1305.wr_en = AESL_inst_myproject.layer2_out_1304_U.if_write & AESL_inst_myproject.layer2_out_1304_U.if_full_n;
    assign fifo_intf_1305.fifo_rd_block = 0;
    assign fifo_intf_1305.fifo_wr_block = 0;
    assign fifo_intf_1305.finish = finish;
    csv_file_dump fifo_csv_dumper_1305;
    csv_file_dump cstatus_csv_dumper_1305;
    df_fifo_monitor fifo_monitor_1305;
    df_fifo_intf fifo_intf_1306(clock,reset);
    assign fifo_intf_1306.rd_en = AESL_inst_myproject.layer2_out_1305_U.if_read & AESL_inst_myproject.layer2_out_1305_U.if_empty_n;
    assign fifo_intf_1306.wr_en = AESL_inst_myproject.layer2_out_1305_U.if_write & AESL_inst_myproject.layer2_out_1305_U.if_full_n;
    assign fifo_intf_1306.fifo_rd_block = 0;
    assign fifo_intf_1306.fifo_wr_block = 0;
    assign fifo_intf_1306.finish = finish;
    csv_file_dump fifo_csv_dumper_1306;
    csv_file_dump cstatus_csv_dumper_1306;
    df_fifo_monitor fifo_monitor_1306;
    df_fifo_intf fifo_intf_1307(clock,reset);
    assign fifo_intf_1307.rd_en = AESL_inst_myproject.layer2_out_1306_U.if_read & AESL_inst_myproject.layer2_out_1306_U.if_empty_n;
    assign fifo_intf_1307.wr_en = AESL_inst_myproject.layer2_out_1306_U.if_write & AESL_inst_myproject.layer2_out_1306_U.if_full_n;
    assign fifo_intf_1307.fifo_rd_block = 0;
    assign fifo_intf_1307.fifo_wr_block = 0;
    assign fifo_intf_1307.finish = finish;
    csv_file_dump fifo_csv_dumper_1307;
    csv_file_dump cstatus_csv_dumper_1307;
    df_fifo_monitor fifo_monitor_1307;
    df_fifo_intf fifo_intf_1308(clock,reset);
    assign fifo_intf_1308.rd_en = AESL_inst_myproject.layer2_out_1307_U.if_read & AESL_inst_myproject.layer2_out_1307_U.if_empty_n;
    assign fifo_intf_1308.wr_en = AESL_inst_myproject.layer2_out_1307_U.if_write & AESL_inst_myproject.layer2_out_1307_U.if_full_n;
    assign fifo_intf_1308.fifo_rd_block = 0;
    assign fifo_intf_1308.fifo_wr_block = 0;
    assign fifo_intf_1308.finish = finish;
    csv_file_dump fifo_csv_dumper_1308;
    csv_file_dump cstatus_csv_dumper_1308;
    df_fifo_monitor fifo_monitor_1308;
    df_fifo_intf fifo_intf_1309(clock,reset);
    assign fifo_intf_1309.rd_en = AESL_inst_myproject.layer2_out_1308_U.if_read & AESL_inst_myproject.layer2_out_1308_U.if_empty_n;
    assign fifo_intf_1309.wr_en = AESL_inst_myproject.layer2_out_1308_U.if_write & AESL_inst_myproject.layer2_out_1308_U.if_full_n;
    assign fifo_intf_1309.fifo_rd_block = 0;
    assign fifo_intf_1309.fifo_wr_block = 0;
    assign fifo_intf_1309.finish = finish;
    csv_file_dump fifo_csv_dumper_1309;
    csv_file_dump cstatus_csv_dumper_1309;
    df_fifo_monitor fifo_monitor_1309;
    df_fifo_intf fifo_intf_1310(clock,reset);
    assign fifo_intf_1310.rd_en = AESL_inst_myproject.layer2_out_1309_U.if_read & AESL_inst_myproject.layer2_out_1309_U.if_empty_n;
    assign fifo_intf_1310.wr_en = AESL_inst_myproject.layer2_out_1309_U.if_write & AESL_inst_myproject.layer2_out_1309_U.if_full_n;
    assign fifo_intf_1310.fifo_rd_block = 0;
    assign fifo_intf_1310.fifo_wr_block = 0;
    assign fifo_intf_1310.finish = finish;
    csv_file_dump fifo_csv_dumper_1310;
    csv_file_dump cstatus_csv_dumper_1310;
    df_fifo_monitor fifo_monitor_1310;
    df_fifo_intf fifo_intf_1311(clock,reset);
    assign fifo_intf_1311.rd_en = AESL_inst_myproject.layer2_out_1310_U.if_read & AESL_inst_myproject.layer2_out_1310_U.if_empty_n;
    assign fifo_intf_1311.wr_en = AESL_inst_myproject.layer2_out_1310_U.if_write & AESL_inst_myproject.layer2_out_1310_U.if_full_n;
    assign fifo_intf_1311.fifo_rd_block = 0;
    assign fifo_intf_1311.fifo_wr_block = 0;
    assign fifo_intf_1311.finish = finish;
    csv_file_dump fifo_csv_dumper_1311;
    csv_file_dump cstatus_csv_dumper_1311;
    df_fifo_monitor fifo_monitor_1311;
    df_fifo_intf fifo_intf_1312(clock,reset);
    assign fifo_intf_1312.rd_en = AESL_inst_myproject.layer2_out_1311_U.if_read & AESL_inst_myproject.layer2_out_1311_U.if_empty_n;
    assign fifo_intf_1312.wr_en = AESL_inst_myproject.layer2_out_1311_U.if_write & AESL_inst_myproject.layer2_out_1311_U.if_full_n;
    assign fifo_intf_1312.fifo_rd_block = 0;
    assign fifo_intf_1312.fifo_wr_block = 0;
    assign fifo_intf_1312.finish = finish;
    csv_file_dump fifo_csv_dumper_1312;
    csv_file_dump cstatus_csv_dumper_1312;
    df_fifo_monitor fifo_monitor_1312;
    df_fifo_intf fifo_intf_1313(clock,reset);
    assign fifo_intf_1313.rd_en = AESL_inst_myproject.layer2_out_1312_U.if_read & AESL_inst_myproject.layer2_out_1312_U.if_empty_n;
    assign fifo_intf_1313.wr_en = AESL_inst_myproject.layer2_out_1312_U.if_write & AESL_inst_myproject.layer2_out_1312_U.if_full_n;
    assign fifo_intf_1313.fifo_rd_block = 0;
    assign fifo_intf_1313.fifo_wr_block = 0;
    assign fifo_intf_1313.finish = finish;
    csv_file_dump fifo_csv_dumper_1313;
    csv_file_dump cstatus_csv_dumper_1313;
    df_fifo_monitor fifo_monitor_1313;
    df_fifo_intf fifo_intf_1314(clock,reset);
    assign fifo_intf_1314.rd_en = AESL_inst_myproject.layer2_out_1313_U.if_read & AESL_inst_myproject.layer2_out_1313_U.if_empty_n;
    assign fifo_intf_1314.wr_en = AESL_inst_myproject.layer2_out_1313_U.if_write & AESL_inst_myproject.layer2_out_1313_U.if_full_n;
    assign fifo_intf_1314.fifo_rd_block = 0;
    assign fifo_intf_1314.fifo_wr_block = 0;
    assign fifo_intf_1314.finish = finish;
    csv_file_dump fifo_csv_dumper_1314;
    csv_file_dump cstatus_csv_dumper_1314;
    df_fifo_monitor fifo_monitor_1314;
    df_fifo_intf fifo_intf_1315(clock,reset);
    assign fifo_intf_1315.rd_en = AESL_inst_myproject.layer2_out_1314_U.if_read & AESL_inst_myproject.layer2_out_1314_U.if_empty_n;
    assign fifo_intf_1315.wr_en = AESL_inst_myproject.layer2_out_1314_U.if_write & AESL_inst_myproject.layer2_out_1314_U.if_full_n;
    assign fifo_intf_1315.fifo_rd_block = 0;
    assign fifo_intf_1315.fifo_wr_block = 0;
    assign fifo_intf_1315.finish = finish;
    csv_file_dump fifo_csv_dumper_1315;
    csv_file_dump cstatus_csv_dumper_1315;
    df_fifo_monitor fifo_monitor_1315;
    df_fifo_intf fifo_intf_1316(clock,reset);
    assign fifo_intf_1316.rd_en = AESL_inst_myproject.layer2_out_1315_U.if_read & AESL_inst_myproject.layer2_out_1315_U.if_empty_n;
    assign fifo_intf_1316.wr_en = AESL_inst_myproject.layer2_out_1315_U.if_write & AESL_inst_myproject.layer2_out_1315_U.if_full_n;
    assign fifo_intf_1316.fifo_rd_block = 0;
    assign fifo_intf_1316.fifo_wr_block = 0;
    assign fifo_intf_1316.finish = finish;
    csv_file_dump fifo_csv_dumper_1316;
    csv_file_dump cstatus_csv_dumper_1316;
    df_fifo_monitor fifo_monitor_1316;
    df_fifo_intf fifo_intf_1317(clock,reset);
    assign fifo_intf_1317.rd_en = AESL_inst_myproject.layer2_out_1316_U.if_read & AESL_inst_myproject.layer2_out_1316_U.if_empty_n;
    assign fifo_intf_1317.wr_en = AESL_inst_myproject.layer2_out_1316_U.if_write & AESL_inst_myproject.layer2_out_1316_U.if_full_n;
    assign fifo_intf_1317.fifo_rd_block = 0;
    assign fifo_intf_1317.fifo_wr_block = 0;
    assign fifo_intf_1317.finish = finish;
    csv_file_dump fifo_csv_dumper_1317;
    csv_file_dump cstatus_csv_dumper_1317;
    df_fifo_monitor fifo_monitor_1317;
    df_fifo_intf fifo_intf_1318(clock,reset);
    assign fifo_intf_1318.rd_en = AESL_inst_myproject.layer2_out_1317_U.if_read & AESL_inst_myproject.layer2_out_1317_U.if_empty_n;
    assign fifo_intf_1318.wr_en = AESL_inst_myproject.layer2_out_1317_U.if_write & AESL_inst_myproject.layer2_out_1317_U.if_full_n;
    assign fifo_intf_1318.fifo_rd_block = 0;
    assign fifo_intf_1318.fifo_wr_block = 0;
    assign fifo_intf_1318.finish = finish;
    csv_file_dump fifo_csv_dumper_1318;
    csv_file_dump cstatus_csv_dumper_1318;
    df_fifo_monitor fifo_monitor_1318;
    df_fifo_intf fifo_intf_1319(clock,reset);
    assign fifo_intf_1319.rd_en = AESL_inst_myproject.layer2_out_1318_U.if_read & AESL_inst_myproject.layer2_out_1318_U.if_empty_n;
    assign fifo_intf_1319.wr_en = AESL_inst_myproject.layer2_out_1318_U.if_write & AESL_inst_myproject.layer2_out_1318_U.if_full_n;
    assign fifo_intf_1319.fifo_rd_block = 0;
    assign fifo_intf_1319.fifo_wr_block = 0;
    assign fifo_intf_1319.finish = finish;
    csv_file_dump fifo_csv_dumper_1319;
    csv_file_dump cstatus_csv_dumper_1319;
    df_fifo_monitor fifo_monitor_1319;
    df_fifo_intf fifo_intf_1320(clock,reset);
    assign fifo_intf_1320.rd_en = AESL_inst_myproject.layer2_out_1319_U.if_read & AESL_inst_myproject.layer2_out_1319_U.if_empty_n;
    assign fifo_intf_1320.wr_en = AESL_inst_myproject.layer2_out_1319_U.if_write & AESL_inst_myproject.layer2_out_1319_U.if_full_n;
    assign fifo_intf_1320.fifo_rd_block = 0;
    assign fifo_intf_1320.fifo_wr_block = 0;
    assign fifo_intf_1320.finish = finish;
    csv_file_dump fifo_csv_dumper_1320;
    csv_file_dump cstatus_csv_dumper_1320;
    df_fifo_monitor fifo_monitor_1320;
    df_fifo_intf fifo_intf_1321(clock,reset);
    assign fifo_intf_1321.rd_en = AESL_inst_myproject.layer2_out_1320_U.if_read & AESL_inst_myproject.layer2_out_1320_U.if_empty_n;
    assign fifo_intf_1321.wr_en = AESL_inst_myproject.layer2_out_1320_U.if_write & AESL_inst_myproject.layer2_out_1320_U.if_full_n;
    assign fifo_intf_1321.fifo_rd_block = 0;
    assign fifo_intf_1321.fifo_wr_block = 0;
    assign fifo_intf_1321.finish = finish;
    csv_file_dump fifo_csv_dumper_1321;
    csv_file_dump cstatus_csv_dumper_1321;
    df_fifo_monitor fifo_monitor_1321;
    df_fifo_intf fifo_intf_1322(clock,reset);
    assign fifo_intf_1322.rd_en = AESL_inst_myproject.layer2_out_1321_U.if_read & AESL_inst_myproject.layer2_out_1321_U.if_empty_n;
    assign fifo_intf_1322.wr_en = AESL_inst_myproject.layer2_out_1321_U.if_write & AESL_inst_myproject.layer2_out_1321_U.if_full_n;
    assign fifo_intf_1322.fifo_rd_block = 0;
    assign fifo_intf_1322.fifo_wr_block = 0;
    assign fifo_intf_1322.finish = finish;
    csv_file_dump fifo_csv_dumper_1322;
    csv_file_dump cstatus_csv_dumper_1322;
    df_fifo_monitor fifo_monitor_1322;
    df_fifo_intf fifo_intf_1323(clock,reset);
    assign fifo_intf_1323.rd_en = AESL_inst_myproject.layer2_out_1322_U.if_read & AESL_inst_myproject.layer2_out_1322_U.if_empty_n;
    assign fifo_intf_1323.wr_en = AESL_inst_myproject.layer2_out_1322_U.if_write & AESL_inst_myproject.layer2_out_1322_U.if_full_n;
    assign fifo_intf_1323.fifo_rd_block = 0;
    assign fifo_intf_1323.fifo_wr_block = 0;
    assign fifo_intf_1323.finish = finish;
    csv_file_dump fifo_csv_dumper_1323;
    csv_file_dump cstatus_csv_dumper_1323;
    df_fifo_monitor fifo_monitor_1323;
    df_fifo_intf fifo_intf_1324(clock,reset);
    assign fifo_intf_1324.rd_en = AESL_inst_myproject.layer2_out_1323_U.if_read & AESL_inst_myproject.layer2_out_1323_U.if_empty_n;
    assign fifo_intf_1324.wr_en = AESL_inst_myproject.layer2_out_1323_U.if_write & AESL_inst_myproject.layer2_out_1323_U.if_full_n;
    assign fifo_intf_1324.fifo_rd_block = 0;
    assign fifo_intf_1324.fifo_wr_block = 0;
    assign fifo_intf_1324.finish = finish;
    csv_file_dump fifo_csv_dumper_1324;
    csv_file_dump cstatus_csv_dumper_1324;
    df_fifo_monitor fifo_monitor_1324;
    df_fifo_intf fifo_intf_1325(clock,reset);
    assign fifo_intf_1325.rd_en = AESL_inst_myproject.layer2_out_1324_U.if_read & AESL_inst_myproject.layer2_out_1324_U.if_empty_n;
    assign fifo_intf_1325.wr_en = AESL_inst_myproject.layer2_out_1324_U.if_write & AESL_inst_myproject.layer2_out_1324_U.if_full_n;
    assign fifo_intf_1325.fifo_rd_block = 0;
    assign fifo_intf_1325.fifo_wr_block = 0;
    assign fifo_intf_1325.finish = finish;
    csv_file_dump fifo_csv_dumper_1325;
    csv_file_dump cstatus_csv_dumper_1325;
    df_fifo_monitor fifo_monitor_1325;
    df_fifo_intf fifo_intf_1326(clock,reset);
    assign fifo_intf_1326.rd_en = AESL_inst_myproject.layer2_out_1325_U.if_read & AESL_inst_myproject.layer2_out_1325_U.if_empty_n;
    assign fifo_intf_1326.wr_en = AESL_inst_myproject.layer2_out_1325_U.if_write & AESL_inst_myproject.layer2_out_1325_U.if_full_n;
    assign fifo_intf_1326.fifo_rd_block = 0;
    assign fifo_intf_1326.fifo_wr_block = 0;
    assign fifo_intf_1326.finish = finish;
    csv_file_dump fifo_csv_dumper_1326;
    csv_file_dump cstatus_csv_dumper_1326;
    df_fifo_monitor fifo_monitor_1326;
    df_fifo_intf fifo_intf_1327(clock,reset);
    assign fifo_intf_1327.rd_en = AESL_inst_myproject.layer2_out_1326_U.if_read & AESL_inst_myproject.layer2_out_1326_U.if_empty_n;
    assign fifo_intf_1327.wr_en = AESL_inst_myproject.layer2_out_1326_U.if_write & AESL_inst_myproject.layer2_out_1326_U.if_full_n;
    assign fifo_intf_1327.fifo_rd_block = 0;
    assign fifo_intf_1327.fifo_wr_block = 0;
    assign fifo_intf_1327.finish = finish;
    csv_file_dump fifo_csv_dumper_1327;
    csv_file_dump cstatus_csv_dumper_1327;
    df_fifo_monitor fifo_monitor_1327;
    df_fifo_intf fifo_intf_1328(clock,reset);
    assign fifo_intf_1328.rd_en = AESL_inst_myproject.layer2_out_1327_U.if_read & AESL_inst_myproject.layer2_out_1327_U.if_empty_n;
    assign fifo_intf_1328.wr_en = AESL_inst_myproject.layer2_out_1327_U.if_write & AESL_inst_myproject.layer2_out_1327_U.if_full_n;
    assign fifo_intf_1328.fifo_rd_block = 0;
    assign fifo_intf_1328.fifo_wr_block = 0;
    assign fifo_intf_1328.finish = finish;
    csv_file_dump fifo_csv_dumper_1328;
    csv_file_dump cstatus_csv_dumper_1328;
    df_fifo_monitor fifo_monitor_1328;
    df_fifo_intf fifo_intf_1329(clock,reset);
    assign fifo_intf_1329.rd_en = AESL_inst_myproject.layer2_out_1328_U.if_read & AESL_inst_myproject.layer2_out_1328_U.if_empty_n;
    assign fifo_intf_1329.wr_en = AESL_inst_myproject.layer2_out_1328_U.if_write & AESL_inst_myproject.layer2_out_1328_U.if_full_n;
    assign fifo_intf_1329.fifo_rd_block = 0;
    assign fifo_intf_1329.fifo_wr_block = 0;
    assign fifo_intf_1329.finish = finish;
    csv_file_dump fifo_csv_dumper_1329;
    csv_file_dump cstatus_csv_dumper_1329;
    df_fifo_monitor fifo_monitor_1329;
    df_fifo_intf fifo_intf_1330(clock,reset);
    assign fifo_intf_1330.rd_en = AESL_inst_myproject.layer2_out_1329_U.if_read & AESL_inst_myproject.layer2_out_1329_U.if_empty_n;
    assign fifo_intf_1330.wr_en = AESL_inst_myproject.layer2_out_1329_U.if_write & AESL_inst_myproject.layer2_out_1329_U.if_full_n;
    assign fifo_intf_1330.fifo_rd_block = 0;
    assign fifo_intf_1330.fifo_wr_block = 0;
    assign fifo_intf_1330.finish = finish;
    csv_file_dump fifo_csv_dumper_1330;
    csv_file_dump cstatus_csv_dumper_1330;
    df_fifo_monitor fifo_monitor_1330;
    df_fifo_intf fifo_intf_1331(clock,reset);
    assign fifo_intf_1331.rd_en = AESL_inst_myproject.layer2_out_1330_U.if_read & AESL_inst_myproject.layer2_out_1330_U.if_empty_n;
    assign fifo_intf_1331.wr_en = AESL_inst_myproject.layer2_out_1330_U.if_write & AESL_inst_myproject.layer2_out_1330_U.if_full_n;
    assign fifo_intf_1331.fifo_rd_block = 0;
    assign fifo_intf_1331.fifo_wr_block = 0;
    assign fifo_intf_1331.finish = finish;
    csv_file_dump fifo_csv_dumper_1331;
    csv_file_dump cstatus_csv_dumper_1331;
    df_fifo_monitor fifo_monitor_1331;
    df_fifo_intf fifo_intf_1332(clock,reset);
    assign fifo_intf_1332.rd_en = AESL_inst_myproject.layer2_out_1331_U.if_read & AESL_inst_myproject.layer2_out_1331_U.if_empty_n;
    assign fifo_intf_1332.wr_en = AESL_inst_myproject.layer2_out_1331_U.if_write & AESL_inst_myproject.layer2_out_1331_U.if_full_n;
    assign fifo_intf_1332.fifo_rd_block = 0;
    assign fifo_intf_1332.fifo_wr_block = 0;
    assign fifo_intf_1332.finish = finish;
    csv_file_dump fifo_csv_dumper_1332;
    csv_file_dump cstatus_csv_dumper_1332;
    df_fifo_monitor fifo_monitor_1332;
    df_fifo_intf fifo_intf_1333(clock,reset);
    assign fifo_intf_1333.rd_en = AESL_inst_myproject.layer2_out_1332_U.if_read & AESL_inst_myproject.layer2_out_1332_U.if_empty_n;
    assign fifo_intf_1333.wr_en = AESL_inst_myproject.layer2_out_1332_U.if_write & AESL_inst_myproject.layer2_out_1332_U.if_full_n;
    assign fifo_intf_1333.fifo_rd_block = 0;
    assign fifo_intf_1333.fifo_wr_block = 0;
    assign fifo_intf_1333.finish = finish;
    csv_file_dump fifo_csv_dumper_1333;
    csv_file_dump cstatus_csv_dumper_1333;
    df_fifo_monitor fifo_monitor_1333;
    df_fifo_intf fifo_intf_1334(clock,reset);
    assign fifo_intf_1334.rd_en = AESL_inst_myproject.layer2_out_1333_U.if_read & AESL_inst_myproject.layer2_out_1333_U.if_empty_n;
    assign fifo_intf_1334.wr_en = AESL_inst_myproject.layer2_out_1333_U.if_write & AESL_inst_myproject.layer2_out_1333_U.if_full_n;
    assign fifo_intf_1334.fifo_rd_block = 0;
    assign fifo_intf_1334.fifo_wr_block = 0;
    assign fifo_intf_1334.finish = finish;
    csv_file_dump fifo_csv_dumper_1334;
    csv_file_dump cstatus_csv_dumper_1334;
    df_fifo_monitor fifo_monitor_1334;
    df_fifo_intf fifo_intf_1335(clock,reset);
    assign fifo_intf_1335.rd_en = AESL_inst_myproject.layer2_out_1334_U.if_read & AESL_inst_myproject.layer2_out_1334_U.if_empty_n;
    assign fifo_intf_1335.wr_en = AESL_inst_myproject.layer2_out_1334_U.if_write & AESL_inst_myproject.layer2_out_1334_U.if_full_n;
    assign fifo_intf_1335.fifo_rd_block = 0;
    assign fifo_intf_1335.fifo_wr_block = 0;
    assign fifo_intf_1335.finish = finish;
    csv_file_dump fifo_csv_dumper_1335;
    csv_file_dump cstatus_csv_dumper_1335;
    df_fifo_monitor fifo_monitor_1335;
    df_fifo_intf fifo_intf_1336(clock,reset);
    assign fifo_intf_1336.rd_en = AESL_inst_myproject.layer2_out_1335_U.if_read & AESL_inst_myproject.layer2_out_1335_U.if_empty_n;
    assign fifo_intf_1336.wr_en = AESL_inst_myproject.layer2_out_1335_U.if_write & AESL_inst_myproject.layer2_out_1335_U.if_full_n;
    assign fifo_intf_1336.fifo_rd_block = 0;
    assign fifo_intf_1336.fifo_wr_block = 0;
    assign fifo_intf_1336.finish = finish;
    csv_file_dump fifo_csv_dumper_1336;
    csv_file_dump cstatus_csv_dumper_1336;
    df_fifo_monitor fifo_monitor_1336;
    df_fifo_intf fifo_intf_1337(clock,reset);
    assign fifo_intf_1337.rd_en = AESL_inst_myproject.layer2_out_1336_U.if_read & AESL_inst_myproject.layer2_out_1336_U.if_empty_n;
    assign fifo_intf_1337.wr_en = AESL_inst_myproject.layer2_out_1336_U.if_write & AESL_inst_myproject.layer2_out_1336_U.if_full_n;
    assign fifo_intf_1337.fifo_rd_block = 0;
    assign fifo_intf_1337.fifo_wr_block = 0;
    assign fifo_intf_1337.finish = finish;
    csv_file_dump fifo_csv_dumper_1337;
    csv_file_dump cstatus_csv_dumper_1337;
    df_fifo_monitor fifo_monitor_1337;
    df_fifo_intf fifo_intf_1338(clock,reset);
    assign fifo_intf_1338.rd_en = AESL_inst_myproject.layer2_out_1337_U.if_read & AESL_inst_myproject.layer2_out_1337_U.if_empty_n;
    assign fifo_intf_1338.wr_en = AESL_inst_myproject.layer2_out_1337_U.if_write & AESL_inst_myproject.layer2_out_1337_U.if_full_n;
    assign fifo_intf_1338.fifo_rd_block = 0;
    assign fifo_intf_1338.fifo_wr_block = 0;
    assign fifo_intf_1338.finish = finish;
    csv_file_dump fifo_csv_dumper_1338;
    csv_file_dump cstatus_csv_dumper_1338;
    df_fifo_monitor fifo_monitor_1338;
    df_fifo_intf fifo_intf_1339(clock,reset);
    assign fifo_intf_1339.rd_en = AESL_inst_myproject.layer2_out_1338_U.if_read & AESL_inst_myproject.layer2_out_1338_U.if_empty_n;
    assign fifo_intf_1339.wr_en = AESL_inst_myproject.layer2_out_1338_U.if_write & AESL_inst_myproject.layer2_out_1338_U.if_full_n;
    assign fifo_intf_1339.fifo_rd_block = 0;
    assign fifo_intf_1339.fifo_wr_block = 0;
    assign fifo_intf_1339.finish = finish;
    csv_file_dump fifo_csv_dumper_1339;
    csv_file_dump cstatus_csv_dumper_1339;
    df_fifo_monitor fifo_monitor_1339;
    df_fifo_intf fifo_intf_1340(clock,reset);
    assign fifo_intf_1340.rd_en = AESL_inst_myproject.layer2_out_1339_U.if_read & AESL_inst_myproject.layer2_out_1339_U.if_empty_n;
    assign fifo_intf_1340.wr_en = AESL_inst_myproject.layer2_out_1339_U.if_write & AESL_inst_myproject.layer2_out_1339_U.if_full_n;
    assign fifo_intf_1340.fifo_rd_block = 0;
    assign fifo_intf_1340.fifo_wr_block = 0;
    assign fifo_intf_1340.finish = finish;
    csv_file_dump fifo_csv_dumper_1340;
    csv_file_dump cstatus_csv_dumper_1340;
    df_fifo_monitor fifo_monitor_1340;
    df_fifo_intf fifo_intf_1341(clock,reset);
    assign fifo_intf_1341.rd_en = AESL_inst_myproject.layer2_out_1340_U.if_read & AESL_inst_myproject.layer2_out_1340_U.if_empty_n;
    assign fifo_intf_1341.wr_en = AESL_inst_myproject.layer2_out_1340_U.if_write & AESL_inst_myproject.layer2_out_1340_U.if_full_n;
    assign fifo_intf_1341.fifo_rd_block = 0;
    assign fifo_intf_1341.fifo_wr_block = 0;
    assign fifo_intf_1341.finish = finish;
    csv_file_dump fifo_csv_dumper_1341;
    csv_file_dump cstatus_csv_dumper_1341;
    df_fifo_monitor fifo_monitor_1341;
    df_fifo_intf fifo_intf_1342(clock,reset);
    assign fifo_intf_1342.rd_en = AESL_inst_myproject.layer2_out_1341_U.if_read & AESL_inst_myproject.layer2_out_1341_U.if_empty_n;
    assign fifo_intf_1342.wr_en = AESL_inst_myproject.layer2_out_1341_U.if_write & AESL_inst_myproject.layer2_out_1341_U.if_full_n;
    assign fifo_intf_1342.fifo_rd_block = 0;
    assign fifo_intf_1342.fifo_wr_block = 0;
    assign fifo_intf_1342.finish = finish;
    csv_file_dump fifo_csv_dumper_1342;
    csv_file_dump cstatus_csv_dumper_1342;
    df_fifo_monitor fifo_monitor_1342;
    df_fifo_intf fifo_intf_1343(clock,reset);
    assign fifo_intf_1343.rd_en = AESL_inst_myproject.layer2_out_1342_U.if_read & AESL_inst_myproject.layer2_out_1342_U.if_empty_n;
    assign fifo_intf_1343.wr_en = AESL_inst_myproject.layer2_out_1342_U.if_write & AESL_inst_myproject.layer2_out_1342_U.if_full_n;
    assign fifo_intf_1343.fifo_rd_block = 0;
    assign fifo_intf_1343.fifo_wr_block = 0;
    assign fifo_intf_1343.finish = finish;
    csv_file_dump fifo_csv_dumper_1343;
    csv_file_dump cstatus_csv_dumper_1343;
    df_fifo_monitor fifo_monitor_1343;
    df_fifo_intf fifo_intf_1344(clock,reset);
    assign fifo_intf_1344.rd_en = AESL_inst_myproject.layer2_out_1343_U.if_read & AESL_inst_myproject.layer2_out_1343_U.if_empty_n;
    assign fifo_intf_1344.wr_en = AESL_inst_myproject.layer2_out_1343_U.if_write & AESL_inst_myproject.layer2_out_1343_U.if_full_n;
    assign fifo_intf_1344.fifo_rd_block = 0;
    assign fifo_intf_1344.fifo_wr_block = 0;
    assign fifo_intf_1344.finish = finish;
    csv_file_dump fifo_csv_dumper_1344;
    csv_file_dump cstatus_csv_dumper_1344;
    df_fifo_monitor fifo_monitor_1344;
    df_fifo_intf fifo_intf_1345(clock,reset);
    assign fifo_intf_1345.rd_en = AESL_inst_myproject.layer2_out_1344_U.if_read & AESL_inst_myproject.layer2_out_1344_U.if_empty_n;
    assign fifo_intf_1345.wr_en = AESL_inst_myproject.layer2_out_1344_U.if_write & AESL_inst_myproject.layer2_out_1344_U.if_full_n;
    assign fifo_intf_1345.fifo_rd_block = 0;
    assign fifo_intf_1345.fifo_wr_block = 0;
    assign fifo_intf_1345.finish = finish;
    csv_file_dump fifo_csv_dumper_1345;
    csv_file_dump cstatus_csv_dumper_1345;
    df_fifo_monitor fifo_monitor_1345;
    df_fifo_intf fifo_intf_1346(clock,reset);
    assign fifo_intf_1346.rd_en = AESL_inst_myproject.layer2_out_1345_U.if_read & AESL_inst_myproject.layer2_out_1345_U.if_empty_n;
    assign fifo_intf_1346.wr_en = AESL_inst_myproject.layer2_out_1345_U.if_write & AESL_inst_myproject.layer2_out_1345_U.if_full_n;
    assign fifo_intf_1346.fifo_rd_block = 0;
    assign fifo_intf_1346.fifo_wr_block = 0;
    assign fifo_intf_1346.finish = finish;
    csv_file_dump fifo_csv_dumper_1346;
    csv_file_dump cstatus_csv_dumper_1346;
    df_fifo_monitor fifo_monitor_1346;
    df_fifo_intf fifo_intf_1347(clock,reset);
    assign fifo_intf_1347.rd_en = AESL_inst_myproject.layer2_out_1346_U.if_read & AESL_inst_myproject.layer2_out_1346_U.if_empty_n;
    assign fifo_intf_1347.wr_en = AESL_inst_myproject.layer2_out_1346_U.if_write & AESL_inst_myproject.layer2_out_1346_U.if_full_n;
    assign fifo_intf_1347.fifo_rd_block = 0;
    assign fifo_intf_1347.fifo_wr_block = 0;
    assign fifo_intf_1347.finish = finish;
    csv_file_dump fifo_csv_dumper_1347;
    csv_file_dump cstatus_csv_dumper_1347;
    df_fifo_monitor fifo_monitor_1347;
    df_fifo_intf fifo_intf_1348(clock,reset);
    assign fifo_intf_1348.rd_en = AESL_inst_myproject.layer2_out_1347_U.if_read & AESL_inst_myproject.layer2_out_1347_U.if_empty_n;
    assign fifo_intf_1348.wr_en = AESL_inst_myproject.layer2_out_1347_U.if_write & AESL_inst_myproject.layer2_out_1347_U.if_full_n;
    assign fifo_intf_1348.fifo_rd_block = 0;
    assign fifo_intf_1348.fifo_wr_block = 0;
    assign fifo_intf_1348.finish = finish;
    csv_file_dump fifo_csv_dumper_1348;
    csv_file_dump cstatus_csv_dumper_1348;
    df_fifo_monitor fifo_monitor_1348;
    df_fifo_intf fifo_intf_1349(clock,reset);
    assign fifo_intf_1349.rd_en = AESL_inst_myproject.layer2_out_1348_U.if_read & AESL_inst_myproject.layer2_out_1348_U.if_empty_n;
    assign fifo_intf_1349.wr_en = AESL_inst_myproject.layer2_out_1348_U.if_write & AESL_inst_myproject.layer2_out_1348_U.if_full_n;
    assign fifo_intf_1349.fifo_rd_block = 0;
    assign fifo_intf_1349.fifo_wr_block = 0;
    assign fifo_intf_1349.finish = finish;
    csv_file_dump fifo_csv_dumper_1349;
    csv_file_dump cstatus_csv_dumper_1349;
    df_fifo_monitor fifo_monitor_1349;
    df_fifo_intf fifo_intf_1350(clock,reset);
    assign fifo_intf_1350.rd_en = AESL_inst_myproject.layer2_out_1349_U.if_read & AESL_inst_myproject.layer2_out_1349_U.if_empty_n;
    assign fifo_intf_1350.wr_en = AESL_inst_myproject.layer2_out_1349_U.if_write & AESL_inst_myproject.layer2_out_1349_U.if_full_n;
    assign fifo_intf_1350.fifo_rd_block = 0;
    assign fifo_intf_1350.fifo_wr_block = 0;
    assign fifo_intf_1350.finish = finish;
    csv_file_dump fifo_csv_dumper_1350;
    csv_file_dump cstatus_csv_dumper_1350;
    df_fifo_monitor fifo_monitor_1350;
    df_fifo_intf fifo_intf_1351(clock,reset);
    assign fifo_intf_1351.rd_en = AESL_inst_myproject.layer2_out_1350_U.if_read & AESL_inst_myproject.layer2_out_1350_U.if_empty_n;
    assign fifo_intf_1351.wr_en = AESL_inst_myproject.layer2_out_1350_U.if_write & AESL_inst_myproject.layer2_out_1350_U.if_full_n;
    assign fifo_intf_1351.fifo_rd_block = 0;
    assign fifo_intf_1351.fifo_wr_block = 0;
    assign fifo_intf_1351.finish = finish;
    csv_file_dump fifo_csv_dumper_1351;
    csv_file_dump cstatus_csv_dumper_1351;
    df_fifo_monitor fifo_monitor_1351;
    df_fifo_intf fifo_intf_1352(clock,reset);
    assign fifo_intf_1352.rd_en = AESL_inst_myproject.layer2_out_1351_U.if_read & AESL_inst_myproject.layer2_out_1351_U.if_empty_n;
    assign fifo_intf_1352.wr_en = AESL_inst_myproject.layer2_out_1351_U.if_write & AESL_inst_myproject.layer2_out_1351_U.if_full_n;
    assign fifo_intf_1352.fifo_rd_block = 0;
    assign fifo_intf_1352.fifo_wr_block = 0;
    assign fifo_intf_1352.finish = finish;
    csv_file_dump fifo_csv_dumper_1352;
    csv_file_dump cstatus_csv_dumper_1352;
    df_fifo_monitor fifo_monitor_1352;
    df_fifo_intf fifo_intf_1353(clock,reset);
    assign fifo_intf_1353.rd_en = AESL_inst_myproject.layer3_out_U.if_read & AESL_inst_myproject.layer3_out_U.if_empty_n;
    assign fifo_intf_1353.wr_en = AESL_inst_myproject.layer3_out_U.if_write & AESL_inst_myproject.layer3_out_U.if_full_n;
    assign fifo_intf_1353.fifo_rd_block = 0;
    assign fifo_intf_1353.fifo_wr_block = 0;
    assign fifo_intf_1353.finish = finish;
    csv_file_dump fifo_csv_dumper_1353;
    csv_file_dump cstatus_csv_dumper_1353;
    df_fifo_monitor fifo_monitor_1353;
    df_fifo_intf fifo_intf_1354(clock,reset);
    assign fifo_intf_1354.rd_en = AESL_inst_myproject.layer3_out_1_U.if_read & AESL_inst_myproject.layer3_out_1_U.if_empty_n;
    assign fifo_intf_1354.wr_en = AESL_inst_myproject.layer3_out_1_U.if_write & AESL_inst_myproject.layer3_out_1_U.if_full_n;
    assign fifo_intf_1354.fifo_rd_block = 0;
    assign fifo_intf_1354.fifo_wr_block = 0;
    assign fifo_intf_1354.finish = finish;
    csv_file_dump fifo_csv_dumper_1354;
    csv_file_dump cstatus_csv_dumper_1354;
    df_fifo_monitor fifo_monitor_1354;
    df_fifo_intf fifo_intf_1355(clock,reset);
    assign fifo_intf_1355.rd_en = AESL_inst_myproject.layer3_out_2_U.if_read & AESL_inst_myproject.layer3_out_2_U.if_empty_n;
    assign fifo_intf_1355.wr_en = AESL_inst_myproject.layer3_out_2_U.if_write & AESL_inst_myproject.layer3_out_2_U.if_full_n;
    assign fifo_intf_1355.fifo_rd_block = 0;
    assign fifo_intf_1355.fifo_wr_block = 0;
    assign fifo_intf_1355.finish = finish;
    csv_file_dump fifo_csv_dumper_1355;
    csv_file_dump cstatus_csv_dumper_1355;
    df_fifo_monitor fifo_monitor_1355;
    df_fifo_intf fifo_intf_1356(clock,reset);
    assign fifo_intf_1356.rd_en = AESL_inst_myproject.layer3_out_3_U.if_read & AESL_inst_myproject.layer3_out_3_U.if_empty_n;
    assign fifo_intf_1356.wr_en = AESL_inst_myproject.layer3_out_3_U.if_write & AESL_inst_myproject.layer3_out_3_U.if_full_n;
    assign fifo_intf_1356.fifo_rd_block = 0;
    assign fifo_intf_1356.fifo_wr_block = 0;
    assign fifo_intf_1356.finish = finish;
    csv_file_dump fifo_csv_dumper_1356;
    csv_file_dump cstatus_csv_dumper_1356;
    df_fifo_monitor fifo_monitor_1356;
    df_fifo_intf fifo_intf_1357(clock,reset);
    assign fifo_intf_1357.rd_en = AESL_inst_myproject.layer3_out_4_U.if_read & AESL_inst_myproject.layer3_out_4_U.if_empty_n;
    assign fifo_intf_1357.wr_en = AESL_inst_myproject.layer3_out_4_U.if_write & AESL_inst_myproject.layer3_out_4_U.if_full_n;
    assign fifo_intf_1357.fifo_rd_block = 0;
    assign fifo_intf_1357.fifo_wr_block = 0;
    assign fifo_intf_1357.finish = finish;
    csv_file_dump fifo_csv_dumper_1357;
    csv_file_dump cstatus_csv_dumper_1357;
    df_fifo_monitor fifo_monitor_1357;
    df_fifo_intf fifo_intf_1358(clock,reset);
    assign fifo_intf_1358.rd_en = AESL_inst_myproject.layer3_out_5_U.if_read & AESL_inst_myproject.layer3_out_5_U.if_empty_n;
    assign fifo_intf_1358.wr_en = AESL_inst_myproject.layer3_out_5_U.if_write & AESL_inst_myproject.layer3_out_5_U.if_full_n;
    assign fifo_intf_1358.fifo_rd_block = 0;
    assign fifo_intf_1358.fifo_wr_block = 0;
    assign fifo_intf_1358.finish = finish;
    csv_file_dump fifo_csv_dumper_1358;
    csv_file_dump cstatus_csv_dumper_1358;
    df_fifo_monitor fifo_monitor_1358;
    df_fifo_intf fifo_intf_1359(clock,reset);
    assign fifo_intf_1359.rd_en = AESL_inst_myproject.layer3_out_6_U.if_read & AESL_inst_myproject.layer3_out_6_U.if_empty_n;
    assign fifo_intf_1359.wr_en = AESL_inst_myproject.layer3_out_6_U.if_write & AESL_inst_myproject.layer3_out_6_U.if_full_n;
    assign fifo_intf_1359.fifo_rd_block = 0;
    assign fifo_intf_1359.fifo_wr_block = 0;
    assign fifo_intf_1359.finish = finish;
    csv_file_dump fifo_csv_dumper_1359;
    csv_file_dump cstatus_csv_dumper_1359;
    df_fifo_monitor fifo_monitor_1359;
    df_fifo_intf fifo_intf_1360(clock,reset);
    assign fifo_intf_1360.rd_en = AESL_inst_myproject.layer3_out_7_U.if_read & AESL_inst_myproject.layer3_out_7_U.if_empty_n;
    assign fifo_intf_1360.wr_en = AESL_inst_myproject.layer3_out_7_U.if_write & AESL_inst_myproject.layer3_out_7_U.if_full_n;
    assign fifo_intf_1360.fifo_rd_block = 0;
    assign fifo_intf_1360.fifo_wr_block = 0;
    assign fifo_intf_1360.finish = finish;
    csv_file_dump fifo_csv_dumper_1360;
    csv_file_dump cstatus_csv_dumper_1360;
    df_fifo_monitor fifo_monitor_1360;
    df_fifo_intf fifo_intf_1361(clock,reset);
    assign fifo_intf_1361.rd_en = AESL_inst_myproject.layer3_out_8_U.if_read & AESL_inst_myproject.layer3_out_8_U.if_empty_n;
    assign fifo_intf_1361.wr_en = AESL_inst_myproject.layer3_out_8_U.if_write & AESL_inst_myproject.layer3_out_8_U.if_full_n;
    assign fifo_intf_1361.fifo_rd_block = 0;
    assign fifo_intf_1361.fifo_wr_block = 0;
    assign fifo_intf_1361.finish = finish;
    csv_file_dump fifo_csv_dumper_1361;
    csv_file_dump cstatus_csv_dumper_1361;
    df_fifo_monitor fifo_monitor_1361;
    df_fifo_intf fifo_intf_1362(clock,reset);
    assign fifo_intf_1362.rd_en = AESL_inst_myproject.layer3_out_9_U.if_read & AESL_inst_myproject.layer3_out_9_U.if_empty_n;
    assign fifo_intf_1362.wr_en = AESL_inst_myproject.layer3_out_9_U.if_write & AESL_inst_myproject.layer3_out_9_U.if_full_n;
    assign fifo_intf_1362.fifo_rd_block = 0;
    assign fifo_intf_1362.fifo_wr_block = 0;
    assign fifo_intf_1362.finish = finish;
    csv_file_dump fifo_csv_dumper_1362;
    csv_file_dump cstatus_csv_dumper_1362;
    df_fifo_monitor fifo_monitor_1362;
    df_fifo_intf fifo_intf_1363(clock,reset);
    assign fifo_intf_1363.rd_en = AESL_inst_myproject.layer3_out_10_U.if_read & AESL_inst_myproject.layer3_out_10_U.if_empty_n;
    assign fifo_intf_1363.wr_en = AESL_inst_myproject.layer3_out_10_U.if_write & AESL_inst_myproject.layer3_out_10_U.if_full_n;
    assign fifo_intf_1363.fifo_rd_block = 0;
    assign fifo_intf_1363.fifo_wr_block = 0;
    assign fifo_intf_1363.finish = finish;
    csv_file_dump fifo_csv_dumper_1363;
    csv_file_dump cstatus_csv_dumper_1363;
    df_fifo_monitor fifo_monitor_1363;
    df_fifo_intf fifo_intf_1364(clock,reset);
    assign fifo_intf_1364.rd_en = AESL_inst_myproject.layer3_out_11_U.if_read & AESL_inst_myproject.layer3_out_11_U.if_empty_n;
    assign fifo_intf_1364.wr_en = AESL_inst_myproject.layer3_out_11_U.if_write & AESL_inst_myproject.layer3_out_11_U.if_full_n;
    assign fifo_intf_1364.fifo_rd_block = 0;
    assign fifo_intf_1364.fifo_wr_block = 0;
    assign fifo_intf_1364.finish = finish;
    csv_file_dump fifo_csv_dumper_1364;
    csv_file_dump cstatus_csv_dumper_1364;
    df_fifo_monitor fifo_monitor_1364;
    df_fifo_intf fifo_intf_1365(clock,reset);
    assign fifo_intf_1365.rd_en = AESL_inst_myproject.layer3_out_12_U.if_read & AESL_inst_myproject.layer3_out_12_U.if_empty_n;
    assign fifo_intf_1365.wr_en = AESL_inst_myproject.layer3_out_12_U.if_write & AESL_inst_myproject.layer3_out_12_U.if_full_n;
    assign fifo_intf_1365.fifo_rd_block = 0;
    assign fifo_intf_1365.fifo_wr_block = 0;
    assign fifo_intf_1365.finish = finish;
    csv_file_dump fifo_csv_dumper_1365;
    csv_file_dump cstatus_csv_dumper_1365;
    df_fifo_monitor fifo_monitor_1365;
    df_fifo_intf fifo_intf_1366(clock,reset);
    assign fifo_intf_1366.rd_en = AESL_inst_myproject.layer3_out_13_U.if_read & AESL_inst_myproject.layer3_out_13_U.if_empty_n;
    assign fifo_intf_1366.wr_en = AESL_inst_myproject.layer3_out_13_U.if_write & AESL_inst_myproject.layer3_out_13_U.if_full_n;
    assign fifo_intf_1366.fifo_rd_block = 0;
    assign fifo_intf_1366.fifo_wr_block = 0;
    assign fifo_intf_1366.finish = finish;
    csv_file_dump fifo_csv_dumper_1366;
    csv_file_dump cstatus_csv_dumper_1366;
    df_fifo_monitor fifo_monitor_1366;
    df_fifo_intf fifo_intf_1367(clock,reset);
    assign fifo_intf_1367.rd_en = AESL_inst_myproject.layer3_out_14_U.if_read & AESL_inst_myproject.layer3_out_14_U.if_empty_n;
    assign fifo_intf_1367.wr_en = AESL_inst_myproject.layer3_out_14_U.if_write & AESL_inst_myproject.layer3_out_14_U.if_full_n;
    assign fifo_intf_1367.fifo_rd_block = 0;
    assign fifo_intf_1367.fifo_wr_block = 0;
    assign fifo_intf_1367.finish = finish;
    csv_file_dump fifo_csv_dumper_1367;
    csv_file_dump cstatus_csv_dumper_1367;
    df_fifo_monitor fifo_monitor_1367;
    df_fifo_intf fifo_intf_1368(clock,reset);
    assign fifo_intf_1368.rd_en = AESL_inst_myproject.layer3_out_15_U.if_read & AESL_inst_myproject.layer3_out_15_U.if_empty_n;
    assign fifo_intf_1368.wr_en = AESL_inst_myproject.layer3_out_15_U.if_write & AESL_inst_myproject.layer3_out_15_U.if_full_n;
    assign fifo_intf_1368.fifo_rd_block = 0;
    assign fifo_intf_1368.fifo_wr_block = 0;
    assign fifo_intf_1368.finish = finish;
    csv_file_dump fifo_csv_dumper_1368;
    csv_file_dump cstatus_csv_dumper_1368;
    df_fifo_monitor fifo_monitor_1368;
    df_fifo_intf fifo_intf_1369(clock,reset);
    assign fifo_intf_1369.rd_en = AESL_inst_myproject.layer3_out_16_U.if_read & AESL_inst_myproject.layer3_out_16_U.if_empty_n;
    assign fifo_intf_1369.wr_en = AESL_inst_myproject.layer3_out_16_U.if_write & AESL_inst_myproject.layer3_out_16_U.if_full_n;
    assign fifo_intf_1369.fifo_rd_block = 0;
    assign fifo_intf_1369.fifo_wr_block = 0;
    assign fifo_intf_1369.finish = finish;
    csv_file_dump fifo_csv_dumper_1369;
    csv_file_dump cstatus_csv_dumper_1369;
    df_fifo_monitor fifo_monitor_1369;
    df_fifo_intf fifo_intf_1370(clock,reset);
    assign fifo_intf_1370.rd_en = AESL_inst_myproject.layer3_out_17_U.if_read & AESL_inst_myproject.layer3_out_17_U.if_empty_n;
    assign fifo_intf_1370.wr_en = AESL_inst_myproject.layer3_out_17_U.if_write & AESL_inst_myproject.layer3_out_17_U.if_full_n;
    assign fifo_intf_1370.fifo_rd_block = 0;
    assign fifo_intf_1370.fifo_wr_block = 0;
    assign fifo_intf_1370.finish = finish;
    csv_file_dump fifo_csv_dumper_1370;
    csv_file_dump cstatus_csv_dumper_1370;
    df_fifo_monitor fifo_monitor_1370;
    df_fifo_intf fifo_intf_1371(clock,reset);
    assign fifo_intf_1371.rd_en = AESL_inst_myproject.layer3_out_18_U.if_read & AESL_inst_myproject.layer3_out_18_U.if_empty_n;
    assign fifo_intf_1371.wr_en = AESL_inst_myproject.layer3_out_18_U.if_write & AESL_inst_myproject.layer3_out_18_U.if_full_n;
    assign fifo_intf_1371.fifo_rd_block = 0;
    assign fifo_intf_1371.fifo_wr_block = 0;
    assign fifo_intf_1371.finish = finish;
    csv_file_dump fifo_csv_dumper_1371;
    csv_file_dump cstatus_csv_dumper_1371;
    df_fifo_monitor fifo_monitor_1371;
    df_fifo_intf fifo_intf_1372(clock,reset);
    assign fifo_intf_1372.rd_en = AESL_inst_myproject.layer3_out_19_U.if_read & AESL_inst_myproject.layer3_out_19_U.if_empty_n;
    assign fifo_intf_1372.wr_en = AESL_inst_myproject.layer3_out_19_U.if_write & AESL_inst_myproject.layer3_out_19_U.if_full_n;
    assign fifo_intf_1372.fifo_rd_block = 0;
    assign fifo_intf_1372.fifo_wr_block = 0;
    assign fifo_intf_1372.finish = finish;
    csv_file_dump fifo_csv_dumper_1372;
    csv_file_dump cstatus_csv_dumper_1372;
    df_fifo_monitor fifo_monitor_1372;
    df_fifo_intf fifo_intf_1373(clock,reset);
    assign fifo_intf_1373.rd_en = AESL_inst_myproject.layer3_out_20_U.if_read & AESL_inst_myproject.layer3_out_20_U.if_empty_n;
    assign fifo_intf_1373.wr_en = AESL_inst_myproject.layer3_out_20_U.if_write & AESL_inst_myproject.layer3_out_20_U.if_full_n;
    assign fifo_intf_1373.fifo_rd_block = 0;
    assign fifo_intf_1373.fifo_wr_block = 0;
    assign fifo_intf_1373.finish = finish;
    csv_file_dump fifo_csv_dumper_1373;
    csv_file_dump cstatus_csv_dumper_1373;
    df_fifo_monitor fifo_monitor_1373;
    df_fifo_intf fifo_intf_1374(clock,reset);
    assign fifo_intf_1374.rd_en = AESL_inst_myproject.layer3_out_21_U.if_read & AESL_inst_myproject.layer3_out_21_U.if_empty_n;
    assign fifo_intf_1374.wr_en = AESL_inst_myproject.layer3_out_21_U.if_write & AESL_inst_myproject.layer3_out_21_U.if_full_n;
    assign fifo_intf_1374.fifo_rd_block = 0;
    assign fifo_intf_1374.fifo_wr_block = 0;
    assign fifo_intf_1374.finish = finish;
    csv_file_dump fifo_csv_dumper_1374;
    csv_file_dump cstatus_csv_dumper_1374;
    df_fifo_monitor fifo_monitor_1374;
    df_fifo_intf fifo_intf_1375(clock,reset);
    assign fifo_intf_1375.rd_en = AESL_inst_myproject.layer3_out_22_U.if_read & AESL_inst_myproject.layer3_out_22_U.if_empty_n;
    assign fifo_intf_1375.wr_en = AESL_inst_myproject.layer3_out_22_U.if_write & AESL_inst_myproject.layer3_out_22_U.if_full_n;
    assign fifo_intf_1375.fifo_rd_block = 0;
    assign fifo_intf_1375.fifo_wr_block = 0;
    assign fifo_intf_1375.finish = finish;
    csv_file_dump fifo_csv_dumper_1375;
    csv_file_dump cstatus_csv_dumper_1375;
    df_fifo_monitor fifo_monitor_1375;
    df_fifo_intf fifo_intf_1376(clock,reset);
    assign fifo_intf_1376.rd_en = AESL_inst_myproject.layer3_out_23_U.if_read & AESL_inst_myproject.layer3_out_23_U.if_empty_n;
    assign fifo_intf_1376.wr_en = AESL_inst_myproject.layer3_out_23_U.if_write & AESL_inst_myproject.layer3_out_23_U.if_full_n;
    assign fifo_intf_1376.fifo_rd_block = 0;
    assign fifo_intf_1376.fifo_wr_block = 0;
    assign fifo_intf_1376.finish = finish;
    csv_file_dump fifo_csv_dumper_1376;
    csv_file_dump cstatus_csv_dumper_1376;
    df_fifo_monitor fifo_monitor_1376;
    df_fifo_intf fifo_intf_1377(clock,reset);
    assign fifo_intf_1377.rd_en = AESL_inst_myproject.layer3_out_24_U.if_read & AESL_inst_myproject.layer3_out_24_U.if_empty_n;
    assign fifo_intf_1377.wr_en = AESL_inst_myproject.layer3_out_24_U.if_write & AESL_inst_myproject.layer3_out_24_U.if_full_n;
    assign fifo_intf_1377.fifo_rd_block = 0;
    assign fifo_intf_1377.fifo_wr_block = 0;
    assign fifo_intf_1377.finish = finish;
    csv_file_dump fifo_csv_dumper_1377;
    csv_file_dump cstatus_csv_dumper_1377;
    df_fifo_monitor fifo_monitor_1377;
    df_fifo_intf fifo_intf_1378(clock,reset);
    assign fifo_intf_1378.rd_en = AESL_inst_myproject.layer3_out_25_U.if_read & AESL_inst_myproject.layer3_out_25_U.if_empty_n;
    assign fifo_intf_1378.wr_en = AESL_inst_myproject.layer3_out_25_U.if_write & AESL_inst_myproject.layer3_out_25_U.if_full_n;
    assign fifo_intf_1378.fifo_rd_block = 0;
    assign fifo_intf_1378.fifo_wr_block = 0;
    assign fifo_intf_1378.finish = finish;
    csv_file_dump fifo_csv_dumper_1378;
    csv_file_dump cstatus_csv_dumper_1378;
    df_fifo_monitor fifo_monitor_1378;
    df_fifo_intf fifo_intf_1379(clock,reset);
    assign fifo_intf_1379.rd_en = AESL_inst_myproject.layer3_out_26_U.if_read & AESL_inst_myproject.layer3_out_26_U.if_empty_n;
    assign fifo_intf_1379.wr_en = AESL_inst_myproject.layer3_out_26_U.if_write & AESL_inst_myproject.layer3_out_26_U.if_full_n;
    assign fifo_intf_1379.fifo_rd_block = 0;
    assign fifo_intf_1379.fifo_wr_block = 0;
    assign fifo_intf_1379.finish = finish;
    csv_file_dump fifo_csv_dumper_1379;
    csv_file_dump cstatus_csv_dumper_1379;
    df_fifo_monitor fifo_monitor_1379;
    df_fifo_intf fifo_intf_1380(clock,reset);
    assign fifo_intf_1380.rd_en = AESL_inst_myproject.layer3_out_27_U.if_read & AESL_inst_myproject.layer3_out_27_U.if_empty_n;
    assign fifo_intf_1380.wr_en = AESL_inst_myproject.layer3_out_27_U.if_write & AESL_inst_myproject.layer3_out_27_U.if_full_n;
    assign fifo_intf_1380.fifo_rd_block = 0;
    assign fifo_intf_1380.fifo_wr_block = 0;
    assign fifo_intf_1380.finish = finish;
    csv_file_dump fifo_csv_dumper_1380;
    csv_file_dump cstatus_csv_dumper_1380;
    df_fifo_monitor fifo_monitor_1380;
    df_fifo_intf fifo_intf_1381(clock,reset);
    assign fifo_intf_1381.rd_en = AESL_inst_myproject.layer3_out_28_U.if_read & AESL_inst_myproject.layer3_out_28_U.if_empty_n;
    assign fifo_intf_1381.wr_en = AESL_inst_myproject.layer3_out_28_U.if_write & AESL_inst_myproject.layer3_out_28_U.if_full_n;
    assign fifo_intf_1381.fifo_rd_block = 0;
    assign fifo_intf_1381.fifo_wr_block = 0;
    assign fifo_intf_1381.finish = finish;
    csv_file_dump fifo_csv_dumper_1381;
    csv_file_dump cstatus_csv_dumper_1381;
    df_fifo_monitor fifo_monitor_1381;
    df_fifo_intf fifo_intf_1382(clock,reset);
    assign fifo_intf_1382.rd_en = AESL_inst_myproject.layer3_out_29_U.if_read & AESL_inst_myproject.layer3_out_29_U.if_empty_n;
    assign fifo_intf_1382.wr_en = AESL_inst_myproject.layer3_out_29_U.if_write & AESL_inst_myproject.layer3_out_29_U.if_full_n;
    assign fifo_intf_1382.fifo_rd_block = 0;
    assign fifo_intf_1382.fifo_wr_block = 0;
    assign fifo_intf_1382.finish = finish;
    csv_file_dump fifo_csv_dumper_1382;
    csv_file_dump cstatus_csv_dumper_1382;
    df_fifo_monitor fifo_monitor_1382;
    df_fifo_intf fifo_intf_1383(clock,reset);
    assign fifo_intf_1383.rd_en = AESL_inst_myproject.layer3_out_30_U.if_read & AESL_inst_myproject.layer3_out_30_U.if_empty_n;
    assign fifo_intf_1383.wr_en = AESL_inst_myproject.layer3_out_30_U.if_write & AESL_inst_myproject.layer3_out_30_U.if_full_n;
    assign fifo_intf_1383.fifo_rd_block = 0;
    assign fifo_intf_1383.fifo_wr_block = 0;
    assign fifo_intf_1383.finish = finish;
    csv_file_dump fifo_csv_dumper_1383;
    csv_file_dump cstatus_csv_dumper_1383;
    df_fifo_monitor fifo_monitor_1383;
    df_fifo_intf fifo_intf_1384(clock,reset);
    assign fifo_intf_1384.rd_en = AESL_inst_myproject.layer3_out_31_U.if_read & AESL_inst_myproject.layer3_out_31_U.if_empty_n;
    assign fifo_intf_1384.wr_en = AESL_inst_myproject.layer3_out_31_U.if_write & AESL_inst_myproject.layer3_out_31_U.if_full_n;
    assign fifo_intf_1384.fifo_rd_block = 0;
    assign fifo_intf_1384.fifo_wr_block = 0;
    assign fifo_intf_1384.finish = finish;
    csv_file_dump fifo_csv_dumper_1384;
    csv_file_dump cstatus_csv_dumper_1384;
    df_fifo_monitor fifo_monitor_1384;
    df_fifo_intf fifo_intf_1385(clock,reset);
    assign fifo_intf_1385.rd_en = AESL_inst_myproject.layer3_out_32_U.if_read & AESL_inst_myproject.layer3_out_32_U.if_empty_n;
    assign fifo_intf_1385.wr_en = AESL_inst_myproject.layer3_out_32_U.if_write & AESL_inst_myproject.layer3_out_32_U.if_full_n;
    assign fifo_intf_1385.fifo_rd_block = 0;
    assign fifo_intf_1385.fifo_wr_block = 0;
    assign fifo_intf_1385.finish = finish;
    csv_file_dump fifo_csv_dumper_1385;
    csv_file_dump cstatus_csv_dumper_1385;
    df_fifo_monitor fifo_monitor_1385;
    df_fifo_intf fifo_intf_1386(clock,reset);
    assign fifo_intf_1386.rd_en = AESL_inst_myproject.layer3_out_33_U.if_read & AESL_inst_myproject.layer3_out_33_U.if_empty_n;
    assign fifo_intf_1386.wr_en = AESL_inst_myproject.layer3_out_33_U.if_write & AESL_inst_myproject.layer3_out_33_U.if_full_n;
    assign fifo_intf_1386.fifo_rd_block = 0;
    assign fifo_intf_1386.fifo_wr_block = 0;
    assign fifo_intf_1386.finish = finish;
    csv_file_dump fifo_csv_dumper_1386;
    csv_file_dump cstatus_csv_dumper_1386;
    df_fifo_monitor fifo_monitor_1386;
    df_fifo_intf fifo_intf_1387(clock,reset);
    assign fifo_intf_1387.rd_en = AESL_inst_myproject.layer3_out_34_U.if_read & AESL_inst_myproject.layer3_out_34_U.if_empty_n;
    assign fifo_intf_1387.wr_en = AESL_inst_myproject.layer3_out_34_U.if_write & AESL_inst_myproject.layer3_out_34_U.if_full_n;
    assign fifo_intf_1387.fifo_rd_block = 0;
    assign fifo_intf_1387.fifo_wr_block = 0;
    assign fifo_intf_1387.finish = finish;
    csv_file_dump fifo_csv_dumper_1387;
    csv_file_dump cstatus_csv_dumper_1387;
    df_fifo_monitor fifo_monitor_1387;
    df_fifo_intf fifo_intf_1388(clock,reset);
    assign fifo_intf_1388.rd_en = AESL_inst_myproject.layer3_out_35_U.if_read & AESL_inst_myproject.layer3_out_35_U.if_empty_n;
    assign fifo_intf_1388.wr_en = AESL_inst_myproject.layer3_out_35_U.if_write & AESL_inst_myproject.layer3_out_35_U.if_full_n;
    assign fifo_intf_1388.fifo_rd_block = 0;
    assign fifo_intf_1388.fifo_wr_block = 0;
    assign fifo_intf_1388.finish = finish;
    csv_file_dump fifo_csv_dumper_1388;
    csv_file_dump cstatus_csv_dumper_1388;
    df_fifo_monitor fifo_monitor_1388;
    df_fifo_intf fifo_intf_1389(clock,reset);
    assign fifo_intf_1389.rd_en = AESL_inst_myproject.layer3_out_36_U.if_read & AESL_inst_myproject.layer3_out_36_U.if_empty_n;
    assign fifo_intf_1389.wr_en = AESL_inst_myproject.layer3_out_36_U.if_write & AESL_inst_myproject.layer3_out_36_U.if_full_n;
    assign fifo_intf_1389.fifo_rd_block = 0;
    assign fifo_intf_1389.fifo_wr_block = 0;
    assign fifo_intf_1389.finish = finish;
    csv_file_dump fifo_csv_dumper_1389;
    csv_file_dump cstatus_csv_dumper_1389;
    df_fifo_monitor fifo_monitor_1389;
    df_fifo_intf fifo_intf_1390(clock,reset);
    assign fifo_intf_1390.rd_en = AESL_inst_myproject.layer3_out_37_U.if_read & AESL_inst_myproject.layer3_out_37_U.if_empty_n;
    assign fifo_intf_1390.wr_en = AESL_inst_myproject.layer3_out_37_U.if_write & AESL_inst_myproject.layer3_out_37_U.if_full_n;
    assign fifo_intf_1390.fifo_rd_block = 0;
    assign fifo_intf_1390.fifo_wr_block = 0;
    assign fifo_intf_1390.finish = finish;
    csv_file_dump fifo_csv_dumper_1390;
    csv_file_dump cstatus_csv_dumper_1390;
    df_fifo_monitor fifo_monitor_1390;
    df_fifo_intf fifo_intf_1391(clock,reset);
    assign fifo_intf_1391.rd_en = AESL_inst_myproject.layer3_out_38_U.if_read & AESL_inst_myproject.layer3_out_38_U.if_empty_n;
    assign fifo_intf_1391.wr_en = AESL_inst_myproject.layer3_out_38_U.if_write & AESL_inst_myproject.layer3_out_38_U.if_full_n;
    assign fifo_intf_1391.fifo_rd_block = 0;
    assign fifo_intf_1391.fifo_wr_block = 0;
    assign fifo_intf_1391.finish = finish;
    csv_file_dump fifo_csv_dumper_1391;
    csv_file_dump cstatus_csv_dumper_1391;
    df_fifo_monitor fifo_monitor_1391;
    df_fifo_intf fifo_intf_1392(clock,reset);
    assign fifo_intf_1392.rd_en = AESL_inst_myproject.layer3_out_39_U.if_read & AESL_inst_myproject.layer3_out_39_U.if_empty_n;
    assign fifo_intf_1392.wr_en = AESL_inst_myproject.layer3_out_39_U.if_write & AESL_inst_myproject.layer3_out_39_U.if_full_n;
    assign fifo_intf_1392.fifo_rd_block = 0;
    assign fifo_intf_1392.fifo_wr_block = 0;
    assign fifo_intf_1392.finish = finish;
    csv_file_dump fifo_csv_dumper_1392;
    csv_file_dump cstatus_csv_dumper_1392;
    df_fifo_monitor fifo_monitor_1392;
    df_fifo_intf fifo_intf_1393(clock,reset);
    assign fifo_intf_1393.rd_en = AESL_inst_myproject.layer3_out_40_U.if_read & AESL_inst_myproject.layer3_out_40_U.if_empty_n;
    assign fifo_intf_1393.wr_en = AESL_inst_myproject.layer3_out_40_U.if_write & AESL_inst_myproject.layer3_out_40_U.if_full_n;
    assign fifo_intf_1393.fifo_rd_block = 0;
    assign fifo_intf_1393.fifo_wr_block = 0;
    assign fifo_intf_1393.finish = finish;
    csv_file_dump fifo_csv_dumper_1393;
    csv_file_dump cstatus_csv_dumper_1393;
    df_fifo_monitor fifo_monitor_1393;
    df_fifo_intf fifo_intf_1394(clock,reset);
    assign fifo_intf_1394.rd_en = AESL_inst_myproject.layer3_out_41_U.if_read & AESL_inst_myproject.layer3_out_41_U.if_empty_n;
    assign fifo_intf_1394.wr_en = AESL_inst_myproject.layer3_out_41_U.if_write & AESL_inst_myproject.layer3_out_41_U.if_full_n;
    assign fifo_intf_1394.fifo_rd_block = 0;
    assign fifo_intf_1394.fifo_wr_block = 0;
    assign fifo_intf_1394.finish = finish;
    csv_file_dump fifo_csv_dumper_1394;
    csv_file_dump cstatus_csv_dumper_1394;
    df_fifo_monitor fifo_monitor_1394;
    df_fifo_intf fifo_intf_1395(clock,reset);
    assign fifo_intf_1395.rd_en = AESL_inst_myproject.layer3_out_42_U.if_read & AESL_inst_myproject.layer3_out_42_U.if_empty_n;
    assign fifo_intf_1395.wr_en = AESL_inst_myproject.layer3_out_42_U.if_write & AESL_inst_myproject.layer3_out_42_U.if_full_n;
    assign fifo_intf_1395.fifo_rd_block = 0;
    assign fifo_intf_1395.fifo_wr_block = 0;
    assign fifo_intf_1395.finish = finish;
    csv_file_dump fifo_csv_dumper_1395;
    csv_file_dump cstatus_csv_dumper_1395;
    df_fifo_monitor fifo_monitor_1395;
    df_fifo_intf fifo_intf_1396(clock,reset);
    assign fifo_intf_1396.rd_en = AESL_inst_myproject.layer3_out_43_U.if_read & AESL_inst_myproject.layer3_out_43_U.if_empty_n;
    assign fifo_intf_1396.wr_en = AESL_inst_myproject.layer3_out_43_U.if_write & AESL_inst_myproject.layer3_out_43_U.if_full_n;
    assign fifo_intf_1396.fifo_rd_block = 0;
    assign fifo_intf_1396.fifo_wr_block = 0;
    assign fifo_intf_1396.finish = finish;
    csv_file_dump fifo_csv_dumper_1396;
    csv_file_dump cstatus_csv_dumper_1396;
    df_fifo_monitor fifo_monitor_1396;
    df_fifo_intf fifo_intf_1397(clock,reset);
    assign fifo_intf_1397.rd_en = AESL_inst_myproject.layer3_out_44_U.if_read & AESL_inst_myproject.layer3_out_44_U.if_empty_n;
    assign fifo_intf_1397.wr_en = AESL_inst_myproject.layer3_out_44_U.if_write & AESL_inst_myproject.layer3_out_44_U.if_full_n;
    assign fifo_intf_1397.fifo_rd_block = 0;
    assign fifo_intf_1397.fifo_wr_block = 0;
    assign fifo_intf_1397.finish = finish;
    csv_file_dump fifo_csv_dumper_1397;
    csv_file_dump cstatus_csv_dumper_1397;
    df_fifo_monitor fifo_monitor_1397;
    df_fifo_intf fifo_intf_1398(clock,reset);
    assign fifo_intf_1398.rd_en = AESL_inst_myproject.layer3_out_45_U.if_read & AESL_inst_myproject.layer3_out_45_U.if_empty_n;
    assign fifo_intf_1398.wr_en = AESL_inst_myproject.layer3_out_45_U.if_write & AESL_inst_myproject.layer3_out_45_U.if_full_n;
    assign fifo_intf_1398.fifo_rd_block = 0;
    assign fifo_intf_1398.fifo_wr_block = 0;
    assign fifo_intf_1398.finish = finish;
    csv_file_dump fifo_csv_dumper_1398;
    csv_file_dump cstatus_csv_dumper_1398;
    df_fifo_monitor fifo_monitor_1398;
    df_fifo_intf fifo_intf_1399(clock,reset);
    assign fifo_intf_1399.rd_en = AESL_inst_myproject.layer3_out_46_U.if_read & AESL_inst_myproject.layer3_out_46_U.if_empty_n;
    assign fifo_intf_1399.wr_en = AESL_inst_myproject.layer3_out_46_U.if_write & AESL_inst_myproject.layer3_out_46_U.if_full_n;
    assign fifo_intf_1399.fifo_rd_block = 0;
    assign fifo_intf_1399.fifo_wr_block = 0;
    assign fifo_intf_1399.finish = finish;
    csv_file_dump fifo_csv_dumper_1399;
    csv_file_dump cstatus_csv_dumper_1399;
    df_fifo_monitor fifo_monitor_1399;
    df_fifo_intf fifo_intf_1400(clock,reset);
    assign fifo_intf_1400.rd_en = AESL_inst_myproject.layer3_out_47_U.if_read & AESL_inst_myproject.layer3_out_47_U.if_empty_n;
    assign fifo_intf_1400.wr_en = AESL_inst_myproject.layer3_out_47_U.if_write & AESL_inst_myproject.layer3_out_47_U.if_full_n;
    assign fifo_intf_1400.fifo_rd_block = 0;
    assign fifo_intf_1400.fifo_wr_block = 0;
    assign fifo_intf_1400.finish = finish;
    csv_file_dump fifo_csv_dumper_1400;
    csv_file_dump cstatus_csv_dumper_1400;
    df_fifo_monitor fifo_monitor_1400;
    df_fifo_intf fifo_intf_1401(clock,reset);
    assign fifo_intf_1401.rd_en = AESL_inst_myproject.layer3_out_48_U.if_read & AESL_inst_myproject.layer3_out_48_U.if_empty_n;
    assign fifo_intf_1401.wr_en = AESL_inst_myproject.layer3_out_48_U.if_write & AESL_inst_myproject.layer3_out_48_U.if_full_n;
    assign fifo_intf_1401.fifo_rd_block = 0;
    assign fifo_intf_1401.fifo_wr_block = 0;
    assign fifo_intf_1401.finish = finish;
    csv_file_dump fifo_csv_dumper_1401;
    csv_file_dump cstatus_csv_dumper_1401;
    df_fifo_monitor fifo_monitor_1401;
    df_fifo_intf fifo_intf_1402(clock,reset);
    assign fifo_intf_1402.rd_en = AESL_inst_myproject.layer3_out_49_U.if_read & AESL_inst_myproject.layer3_out_49_U.if_empty_n;
    assign fifo_intf_1402.wr_en = AESL_inst_myproject.layer3_out_49_U.if_write & AESL_inst_myproject.layer3_out_49_U.if_full_n;
    assign fifo_intf_1402.fifo_rd_block = 0;
    assign fifo_intf_1402.fifo_wr_block = 0;
    assign fifo_intf_1402.finish = finish;
    csv_file_dump fifo_csv_dumper_1402;
    csv_file_dump cstatus_csv_dumper_1402;
    df_fifo_monitor fifo_monitor_1402;
    df_fifo_intf fifo_intf_1403(clock,reset);
    assign fifo_intf_1403.rd_en = AESL_inst_myproject.layer3_out_50_U.if_read & AESL_inst_myproject.layer3_out_50_U.if_empty_n;
    assign fifo_intf_1403.wr_en = AESL_inst_myproject.layer3_out_50_U.if_write & AESL_inst_myproject.layer3_out_50_U.if_full_n;
    assign fifo_intf_1403.fifo_rd_block = 0;
    assign fifo_intf_1403.fifo_wr_block = 0;
    assign fifo_intf_1403.finish = finish;
    csv_file_dump fifo_csv_dumper_1403;
    csv_file_dump cstatus_csv_dumper_1403;
    df_fifo_monitor fifo_monitor_1403;
    df_fifo_intf fifo_intf_1404(clock,reset);
    assign fifo_intf_1404.rd_en = AESL_inst_myproject.layer3_out_51_U.if_read & AESL_inst_myproject.layer3_out_51_U.if_empty_n;
    assign fifo_intf_1404.wr_en = AESL_inst_myproject.layer3_out_51_U.if_write & AESL_inst_myproject.layer3_out_51_U.if_full_n;
    assign fifo_intf_1404.fifo_rd_block = 0;
    assign fifo_intf_1404.fifo_wr_block = 0;
    assign fifo_intf_1404.finish = finish;
    csv_file_dump fifo_csv_dumper_1404;
    csv_file_dump cstatus_csv_dumper_1404;
    df_fifo_monitor fifo_monitor_1404;
    df_fifo_intf fifo_intf_1405(clock,reset);
    assign fifo_intf_1405.rd_en = AESL_inst_myproject.layer3_out_52_U.if_read & AESL_inst_myproject.layer3_out_52_U.if_empty_n;
    assign fifo_intf_1405.wr_en = AESL_inst_myproject.layer3_out_52_U.if_write & AESL_inst_myproject.layer3_out_52_U.if_full_n;
    assign fifo_intf_1405.fifo_rd_block = 0;
    assign fifo_intf_1405.fifo_wr_block = 0;
    assign fifo_intf_1405.finish = finish;
    csv_file_dump fifo_csv_dumper_1405;
    csv_file_dump cstatus_csv_dumper_1405;
    df_fifo_monitor fifo_monitor_1405;
    df_fifo_intf fifo_intf_1406(clock,reset);
    assign fifo_intf_1406.rd_en = AESL_inst_myproject.layer3_out_53_U.if_read & AESL_inst_myproject.layer3_out_53_U.if_empty_n;
    assign fifo_intf_1406.wr_en = AESL_inst_myproject.layer3_out_53_U.if_write & AESL_inst_myproject.layer3_out_53_U.if_full_n;
    assign fifo_intf_1406.fifo_rd_block = 0;
    assign fifo_intf_1406.fifo_wr_block = 0;
    assign fifo_intf_1406.finish = finish;
    csv_file_dump fifo_csv_dumper_1406;
    csv_file_dump cstatus_csv_dumper_1406;
    df_fifo_monitor fifo_monitor_1406;
    df_fifo_intf fifo_intf_1407(clock,reset);
    assign fifo_intf_1407.rd_en = AESL_inst_myproject.layer3_out_54_U.if_read & AESL_inst_myproject.layer3_out_54_U.if_empty_n;
    assign fifo_intf_1407.wr_en = AESL_inst_myproject.layer3_out_54_U.if_write & AESL_inst_myproject.layer3_out_54_U.if_full_n;
    assign fifo_intf_1407.fifo_rd_block = 0;
    assign fifo_intf_1407.fifo_wr_block = 0;
    assign fifo_intf_1407.finish = finish;
    csv_file_dump fifo_csv_dumper_1407;
    csv_file_dump cstatus_csv_dumper_1407;
    df_fifo_monitor fifo_monitor_1407;
    df_fifo_intf fifo_intf_1408(clock,reset);
    assign fifo_intf_1408.rd_en = AESL_inst_myproject.layer3_out_55_U.if_read & AESL_inst_myproject.layer3_out_55_U.if_empty_n;
    assign fifo_intf_1408.wr_en = AESL_inst_myproject.layer3_out_55_U.if_write & AESL_inst_myproject.layer3_out_55_U.if_full_n;
    assign fifo_intf_1408.fifo_rd_block = 0;
    assign fifo_intf_1408.fifo_wr_block = 0;
    assign fifo_intf_1408.finish = finish;
    csv_file_dump fifo_csv_dumper_1408;
    csv_file_dump cstatus_csv_dumper_1408;
    df_fifo_monitor fifo_monitor_1408;
    df_fifo_intf fifo_intf_1409(clock,reset);
    assign fifo_intf_1409.rd_en = AESL_inst_myproject.layer3_out_56_U.if_read & AESL_inst_myproject.layer3_out_56_U.if_empty_n;
    assign fifo_intf_1409.wr_en = AESL_inst_myproject.layer3_out_56_U.if_write & AESL_inst_myproject.layer3_out_56_U.if_full_n;
    assign fifo_intf_1409.fifo_rd_block = 0;
    assign fifo_intf_1409.fifo_wr_block = 0;
    assign fifo_intf_1409.finish = finish;
    csv_file_dump fifo_csv_dumper_1409;
    csv_file_dump cstatus_csv_dumper_1409;
    df_fifo_monitor fifo_monitor_1409;
    df_fifo_intf fifo_intf_1410(clock,reset);
    assign fifo_intf_1410.rd_en = AESL_inst_myproject.layer3_out_57_U.if_read & AESL_inst_myproject.layer3_out_57_U.if_empty_n;
    assign fifo_intf_1410.wr_en = AESL_inst_myproject.layer3_out_57_U.if_write & AESL_inst_myproject.layer3_out_57_U.if_full_n;
    assign fifo_intf_1410.fifo_rd_block = 0;
    assign fifo_intf_1410.fifo_wr_block = 0;
    assign fifo_intf_1410.finish = finish;
    csv_file_dump fifo_csv_dumper_1410;
    csv_file_dump cstatus_csv_dumper_1410;
    df_fifo_monitor fifo_monitor_1410;
    df_fifo_intf fifo_intf_1411(clock,reset);
    assign fifo_intf_1411.rd_en = AESL_inst_myproject.layer3_out_58_U.if_read & AESL_inst_myproject.layer3_out_58_U.if_empty_n;
    assign fifo_intf_1411.wr_en = AESL_inst_myproject.layer3_out_58_U.if_write & AESL_inst_myproject.layer3_out_58_U.if_full_n;
    assign fifo_intf_1411.fifo_rd_block = 0;
    assign fifo_intf_1411.fifo_wr_block = 0;
    assign fifo_intf_1411.finish = finish;
    csv_file_dump fifo_csv_dumper_1411;
    csv_file_dump cstatus_csv_dumper_1411;
    df_fifo_monitor fifo_monitor_1411;
    df_fifo_intf fifo_intf_1412(clock,reset);
    assign fifo_intf_1412.rd_en = AESL_inst_myproject.layer3_out_59_U.if_read & AESL_inst_myproject.layer3_out_59_U.if_empty_n;
    assign fifo_intf_1412.wr_en = AESL_inst_myproject.layer3_out_59_U.if_write & AESL_inst_myproject.layer3_out_59_U.if_full_n;
    assign fifo_intf_1412.fifo_rd_block = 0;
    assign fifo_intf_1412.fifo_wr_block = 0;
    assign fifo_intf_1412.finish = finish;
    csv_file_dump fifo_csv_dumper_1412;
    csv_file_dump cstatus_csv_dumper_1412;
    df_fifo_monitor fifo_monitor_1412;
    df_fifo_intf fifo_intf_1413(clock,reset);
    assign fifo_intf_1413.rd_en = AESL_inst_myproject.layer3_out_60_U.if_read & AESL_inst_myproject.layer3_out_60_U.if_empty_n;
    assign fifo_intf_1413.wr_en = AESL_inst_myproject.layer3_out_60_U.if_write & AESL_inst_myproject.layer3_out_60_U.if_full_n;
    assign fifo_intf_1413.fifo_rd_block = 0;
    assign fifo_intf_1413.fifo_wr_block = 0;
    assign fifo_intf_1413.finish = finish;
    csv_file_dump fifo_csv_dumper_1413;
    csv_file_dump cstatus_csv_dumper_1413;
    df_fifo_monitor fifo_monitor_1413;
    df_fifo_intf fifo_intf_1414(clock,reset);
    assign fifo_intf_1414.rd_en = AESL_inst_myproject.layer3_out_61_U.if_read & AESL_inst_myproject.layer3_out_61_U.if_empty_n;
    assign fifo_intf_1414.wr_en = AESL_inst_myproject.layer3_out_61_U.if_write & AESL_inst_myproject.layer3_out_61_U.if_full_n;
    assign fifo_intf_1414.fifo_rd_block = 0;
    assign fifo_intf_1414.fifo_wr_block = 0;
    assign fifo_intf_1414.finish = finish;
    csv_file_dump fifo_csv_dumper_1414;
    csv_file_dump cstatus_csv_dumper_1414;
    df_fifo_monitor fifo_monitor_1414;
    df_fifo_intf fifo_intf_1415(clock,reset);
    assign fifo_intf_1415.rd_en = AESL_inst_myproject.layer3_out_62_U.if_read & AESL_inst_myproject.layer3_out_62_U.if_empty_n;
    assign fifo_intf_1415.wr_en = AESL_inst_myproject.layer3_out_62_U.if_write & AESL_inst_myproject.layer3_out_62_U.if_full_n;
    assign fifo_intf_1415.fifo_rd_block = 0;
    assign fifo_intf_1415.fifo_wr_block = 0;
    assign fifo_intf_1415.finish = finish;
    csv_file_dump fifo_csv_dumper_1415;
    csv_file_dump cstatus_csv_dumper_1415;
    df_fifo_monitor fifo_monitor_1415;
    df_fifo_intf fifo_intf_1416(clock,reset);
    assign fifo_intf_1416.rd_en = AESL_inst_myproject.layer3_out_63_U.if_read & AESL_inst_myproject.layer3_out_63_U.if_empty_n;
    assign fifo_intf_1416.wr_en = AESL_inst_myproject.layer3_out_63_U.if_write & AESL_inst_myproject.layer3_out_63_U.if_full_n;
    assign fifo_intf_1416.fifo_rd_block = 0;
    assign fifo_intf_1416.fifo_wr_block = 0;
    assign fifo_intf_1416.finish = finish;
    csv_file_dump fifo_csv_dumper_1416;
    csv_file_dump cstatus_csv_dumper_1416;
    df_fifo_monitor fifo_monitor_1416;
    df_fifo_intf fifo_intf_1417(clock,reset);
    assign fifo_intf_1417.rd_en = AESL_inst_myproject.layer3_out_64_U.if_read & AESL_inst_myproject.layer3_out_64_U.if_empty_n;
    assign fifo_intf_1417.wr_en = AESL_inst_myproject.layer3_out_64_U.if_write & AESL_inst_myproject.layer3_out_64_U.if_full_n;
    assign fifo_intf_1417.fifo_rd_block = 0;
    assign fifo_intf_1417.fifo_wr_block = 0;
    assign fifo_intf_1417.finish = finish;
    csv_file_dump fifo_csv_dumper_1417;
    csv_file_dump cstatus_csv_dumper_1417;
    df_fifo_monitor fifo_monitor_1417;
    df_fifo_intf fifo_intf_1418(clock,reset);
    assign fifo_intf_1418.rd_en = AESL_inst_myproject.layer3_out_65_U.if_read & AESL_inst_myproject.layer3_out_65_U.if_empty_n;
    assign fifo_intf_1418.wr_en = AESL_inst_myproject.layer3_out_65_U.if_write & AESL_inst_myproject.layer3_out_65_U.if_full_n;
    assign fifo_intf_1418.fifo_rd_block = 0;
    assign fifo_intf_1418.fifo_wr_block = 0;
    assign fifo_intf_1418.finish = finish;
    csv_file_dump fifo_csv_dumper_1418;
    csv_file_dump cstatus_csv_dumper_1418;
    df_fifo_monitor fifo_monitor_1418;
    df_fifo_intf fifo_intf_1419(clock,reset);
    assign fifo_intf_1419.rd_en = AESL_inst_myproject.layer3_out_66_U.if_read & AESL_inst_myproject.layer3_out_66_U.if_empty_n;
    assign fifo_intf_1419.wr_en = AESL_inst_myproject.layer3_out_66_U.if_write & AESL_inst_myproject.layer3_out_66_U.if_full_n;
    assign fifo_intf_1419.fifo_rd_block = 0;
    assign fifo_intf_1419.fifo_wr_block = 0;
    assign fifo_intf_1419.finish = finish;
    csv_file_dump fifo_csv_dumper_1419;
    csv_file_dump cstatus_csv_dumper_1419;
    df_fifo_monitor fifo_monitor_1419;
    df_fifo_intf fifo_intf_1420(clock,reset);
    assign fifo_intf_1420.rd_en = AESL_inst_myproject.layer3_out_67_U.if_read & AESL_inst_myproject.layer3_out_67_U.if_empty_n;
    assign fifo_intf_1420.wr_en = AESL_inst_myproject.layer3_out_67_U.if_write & AESL_inst_myproject.layer3_out_67_U.if_full_n;
    assign fifo_intf_1420.fifo_rd_block = 0;
    assign fifo_intf_1420.fifo_wr_block = 0;
    assign fifo_intf_1420.finish = finish;
    csv_file_dump fifo_csv_dumper_1420;
    csv_file_dump cstatus_csv_dumper_1420;
    df_fifo_monitor fifo_monitor_1420;
    df_fifo_intf fifo_intf_1421(clock,reset);
    assign fifo_intf_1421.rd_en = AESL_inst_myproject.layer3_out_68_U.if_read & AESL_inst_myproject.layer3_out_68_U.if_empty_n;
    assign fifo_intf_1421.wr_en = AESL_inst_myproject.layer3_out_68_U.if_write & AESL_inst_myproject.layer3_out_68_U.if_full_n;
    assign fifo_intf_1421.fifo_rd_block = 0;
    assign fifo_intf_1421.fifo_wr_block = 0;
    assign fifo_intf_1421.finish = finish;
    csv_file_dump fifo_csv_dumper_1421;
    csv_file_dump cstatus_csv_dumper_1421;
    df_fifo_monitor fifo_monitor_1421;
    df_fifo_intf fifo_intf_1422(clock,reset);
    assign fifo_intf_1422.rd_en = AESL_inst_myproject.layer3_out_69_U.if_read & AESL_inst_myproject.layer3_out_69_U.if_empty_n;
    assign fifo_intf_1422.wr_en = AESL_inst_myproject.layer3_out_69_U.if_write & AESL_inst_myproject.layer3_out_69_U.if_full_n;
    assign fifo_intf_1422.fifo_rd_block = 0;
    assign fifo_intf_1422.fifo_wr_block = 0;
    assign fifo_intf_1422.finish = finish;
    csv_file_dump fifo_csv_dumper_1422;
    csv_file_dump cstatus_csv_dumper_1422;
    df_fifo_monitor fifo_monitor_1422;
    df_fifo_intf fifo_intf_1423(clock,reset);
    assign fifo_intf_1423.rd_en = AESL_inst_myproject.layer3_out_70_U.if_read & AESL_inst_myproject.layer3_out_70_U.if_empty_n;
    assign fifo_intf_1423.wr_en = AESL_inst_myproject.layer3_out_70_U.if_write & AESL_inst_myproject.layer3_out_70_U.if_full_n;
    assign fifo_intf_1423.fifo_rd_block = 0;
    assign fifo_intf_1423.fifo_wr_block = 0;
    assign fifo_intf_1423.finish = finish;
    csv_file_dump fifo_csv_dumper_1423;
    csv_file_dump cstatus_csv_dumper_1423;
    df_fifo_monitor fifo_monitor_1423;
    df_fifo_intf fifo_intf_1424(clock,reset);
    assign fifo_intf_1424.rd_en = AESL_inst_myproject.layer3_out_71_U.if_read & AESL_inst_myproject.layer3_out_71_U.if_empty_n;
    assign fifo_intf_1424.wr_en = AESL_inst_myproject.layer3_out_71_U.if_write & AESL_inst_myproject.layer3_out_71_U.if_full_n;
    assign fifo_intf_1424.fifo_rd_block = 0;
    assign fifo_intf_1424.fifo_wr_block = 0;
    assign fifo_intf_1424.finish = finish;
    csv_file_dump fifo_csv_dumper_1424;
    csv_file_dump cstatus_csv_dumper_1424;
    df_fifo_monitor fifo_monitor_1424;
    df_fifo_intf fifo_intf_1425(clock,reset);
    assign fifo_intf_1425.rd_en = AESL_inst_myproject.layer3_out_72_U.if_read & AESL_inst_myproject.layer3_out_72_U.if_empty_n;
    assign fifo_intf_1425.wr_en = AESL_inst_myproject.layer3_out_72_U.if_write & AESL_inst_myproject.layer3_out_72_U.if_full_n;
    assign fifo_intf_1425.fifo_rd_block = 0;
    assign fifo_intf_1425.fifo_wr_block = 0;
    assign fifo_intf_1425.finish = finish;
    csv_file_dump fifo_csv_dumper_1425;
    csv_file_dump cstatus_csv_dumper_1425;
    df_fifo_monitor fifo_monitor_1425;
    df_fifo_intf fifo_intf_1426(clock,reset);
    assign fifo_intf_1426.rd_en = AESL_inst_myproject.layer3_out_73_U.if_read & AESL_inst_myproject.layer3_out_73_U.if_empty_n;
    assign fifo_intf_1426.wr_en = AESL_inst_myproject.layer3_out_73_U.if_write & AESL_inst_myproject.layer3_out_73_U.if_full_n;
    assign fifo_intf_1426.fifo_rd_block = 0;
    assign fifo_intf_1426.fifo_wr_block = 0;
    assign fifo_intf_1426.finish = finish;
    csv_file_dump fifo_csv_dumper_1426;
    csv_file_dump cstatus_csv_dumper_1426;
    df_fifo_monitor fifo_monitor_1426;
    df_fifo_intf fifo_intf_1427(clock,reset);
    assign fifo_intf_1427.rd_en = AESL_inst_myproject.layer3_out_74_U.if_read & AESL_inst_myproject.layer3_out_74_U.if_empty_n;
    assign fifo_intf_1427.wr_en = AESL_inst_myproject.layer3_out_74_U.if_write & AESL_inst_myproject.layer3_out_74_U.if_full_n;
    assign fifo_intf_1427.fifo_rd_block = 0;
    assign fifo_intf_1427.fifo_wr_block = 0;
    assign fifo_intf_1427.finish = finish;
    csv_file_dump fifo_csv_dumper_1427;
    csv_file_dump cstatus_csv_dumper_1427;
    df_fifo_monitor fifo_monitor_1427;
    df_fifo_intf fifo_intf_1428(clock,reset);
    assign fifo_intf_1428.rd_en = AESL_inst_myproject.layer3_out_75_U.if_read & AESL_inst_myproject.layer3_out_75_U.if_empty_n;
    assign fifo_intf_1428.wr_en = AESL_inst_myproject.layer3_out_75_U.if_write & AESL_inst_myproject.layer3_out_75_U.if_full_n;
    assign fifo_intf_1428.fifo_rd_block = 0;
    assign fifo_intf_1428.fifo_wr_block = 0;
    assign fifo_intf_1428.finish = finish;
    csv_file_dump fifo_csv_dumper_1428;
    csv_file_dump cstatus_csv_dumper_1428;
    df_fifo_monitor fifo_monitor_1428;
    df_fifo_intf fifo_intf_1429(clock,reset);
    assign fifo_intf_1429.rd_en = AESL_inst_myproject.layer3_out_76_U.if_read & AESL_inst_myproject.layer3_out_76_U.if_empty_n;
    assign fifo_intf_1429.wr_en = AESL_inst_myproject.layer3_out_76_U.if_write & AESL_inst_myproject.layer3_out_76_U.if_full_n;
    assign fifo_intf_1429.fifo_rd_block = 0;
    assign fifo_intf_1429.fifo_wr_block = 0;
    assign fifo_intf_1429.finish = finish;
    csv_file_dump fifo_csv_dumper_1429;
    csv_file_dump cstatus_csv_dumper_1429;
    df_fifo_monitor fifo_monitor_1429;
    df_fifo_intf fifo_intf_1430(clock,reset);
    assign fifo_intf_1430.rd_en = AESL_inst_myproject.layer3_out_77_U.if_read & AESL_inst_myproject.layer3_out_77_U.if_empty_n;
    assign fifo_intf_1430.wr_en = AESL_inst_myproject.layer3_out_77_U.if_write & AESL_inst_myproject.layer3_out_77_U.if_full_n;
    assign fifo_intf_1430.fifo_rd_block = 0;
    assign fifo_intf_1430.fifo_wr_block = 0;
    assign fifo_intf_1430.finish = finish;
    csv_file_dump fifo_csv_dumper_1430;
    csv_file_dump cstatus_csv_dumper_1430;
    df_fifo_monitor fifo_monitor_1430;
    df_fifo_intf fifo_intf_1431(clock,reset);
    assign fifo_intf_1431.rd_en = AESL_inst_myproject.layer3_out_78_U.if_read & AESL_inst_myproject.layer3_out_78_U.if_empty_n;
    assign fifo_intf_1431.wr_en = AESL_inst_myproject.layer3_out_78_U.if_write & AESL_inst_myproject.layer3_out_78_U.if_full_n;
    assign fifo_intf_1431.fifo_rd_block = 0;
    assign fifo_intf_1431.fifo_wr_block = 0;
    assign fifo_intf_1431.finish = finish;
    csv_file_dump fifo_csv_dumper_1431;
    csv_file_dump cstatus_csv_dumper_1431;
    df_fifo_monitor fifo_monitor_1431;
    df_fifo_intf fifo_intf_1432(clock,reset);
    assign fifo_intf_1432.rd_en = AESL_inst_myproject.layer3_out_79_U.if_read & AESL_inst_myproject.layer3_out_79_U.if_empty_n;
    assign fifo_intf_1432.wr_en = AESL_inst_myproject.layer3_out_79_U.if_write & AESL_inst_myproject.layer3_out_79_U.if_full_n;
    assign fifo_intf_1432.fifo_rd_block = 0;
    assign fifo_intf_1432.fifo_wr_block = 0;
    assign fifo_intf_1432.finish = finish;
    csv_file_dump fifo_csv_dumper_1432;
    csv_file_dump cstatus_csv_dumper_1432;
    df_fifo_monitor fifo_monitor_1432;
    df_fifo_intf fifo_intf_1433(clock,reset);
    assign fifo_intf_1433.rd_en = AESL_inst_myproject.layer3_out_80_U.if_read & AESL_inst_myproject.layer3_out_80_U.if_empty_n;
    assign fifo_intf_1433.wr_en = AESL_inst_myproject.layer3_out_80_U.if_write & AESL_inst_myproject.layer3_out_80_U.if_full_n;
    assign fifo_intf_1433.fifo_rd_block = 0;
    assign fifo_intf_1433.fifo_wr_block = 0;
    assign fifo_intf_1433.finish = finish;
    csv_file_dump fifo_csv_dumper_1433;
    csv_file_dump cstatus_csv_dumper_1433;
    df_fifo_monitor fifo_monitor_1433;
    df_fifo_intf fifo_intf_1434(clock,reset);
    assign fifo_intf_1434.rd_en = AESL_inst_myproject.layer3_out_81_U.if_read & AESL_inst_myproject.layer3_out_81_U.if_empty_n;
    assign fifo_intf_1434.wr_en = AESL_inst_myproject.layer3_out_81_U.if_write & AESL_inst_myproject.layer3_out_81_U.if_full_n;
    assign fifo_intf_1434.fifo_rd_block = 0;
    assign fifo_intf_1434.fifo_wr_block = 0;
    assign fifo_intf_1434.finish = finish;
    csv_file_dump fifo_csv_dumper_1434;
    csv_file_dump cstatus_csv_dumper_1434;
    df_fifo_monitor fifo_monitor_1434;
    df_fifo_intf fifo_intf_1435(clock,reset);
    assign fifo_intf_1435.rd_en = AESL_inst_myproject.layer3_out_82_U.if_read & AESL_inst_myproject.layer3_out_82_U.if_empty_n;
    assign fifo_intf_1435.wr_en = AESL_inst_myproject.layer3_out_82_U.if_write & AESL_inst_myproject.layer3_out_82_U.if_full_n;
    assign fifo_intf_1435.fifo_rd_block = 0;
    assign fifo_intf_1435.fifo_wr_block = 0;
    assign fifo_intf_1435.finish = finish;
    csv_file_dump fifo_csv_dumper_1435;
    csv_file_dump cstatus_csv_dumper_1435;
    df_fifo_monitor fifo_monitor_1435;
    df_fifo_intf fifo_intf_1436(clock,reset);
    assign fifo_intf_1436.rd_en = AESL_inst_myproject.layer3_out_83_U.if_read & AESL_inst_myproject.layer3_out_83_U.if_empty_n;
    assign fifo_intf_1436.wr_en = AESL_inst_myproject.layer3_out_83_U.if_write & AESL_inst_myproject.layer3_out_83_U.if_full_n;
    assign fifo_intf_1436.fifo_rd_block = 0;
    assign fifo_intf_1436.fifo_wr_block = 0;
    assign fifo_intf_1436.finish = finish;
    csv_file_dump fifo_csv_dumper_1436;
    csv_file_dump cstatus_csv_dumper_1436;
    df_fifo_monitor fifo_monitor_1436;
    df_fifo_intf fifo_intf_1437(clock,reset);
    assign fifo_intf_1437.rd_en = AESL_inst_myproject.layer3_out_84_U.if_read & AESL_inst_myproject.layer3_out_84_U.if_empty_n;
    assign fifo_intf_1437.wr_en = AESL_inst_myproject.layer3_out_84_U.if_write & AESL_inst_myproject.layer3_out_84_U.if_full_n;
    assign fifo_intf_1437.fifo_rd_block = 0;
    assign fifo_intf_1437.fifo_wr_block = 0;
    assign fifo_intf_1437.finish = finish;
    csv_file_dump fifo_csv_dumper_1437;
    csv_file_dump cstatus_csv_dumper_1437;
    df_fifo_monitor fifo_monitor_1437;
    df_fifo_intf fifo_intf_1438(clock,reset);
    assign fifo_intf_1438.rd_en = AESL_inst_myproject.layer3_out_85_U.if_read & AESL_inst_myproject.layer3_out_85_U.if_empty_n;
    assign fifo_intf_1438.wr_en = AESL_inst_myproject.layer3_out_85_U.if_write & AESL_inst_myproject.layer3_out_85_U.if_full_n;
    assign fifo_intf_1438.fifo_rd_block = 0;
    assign fifo_intf_1438.fifo_wr_block = 0;
    assign fifo_intf_1438.finish = finish;
    csv_file_dump fifo_csv_dumper_1438;
    csv_file_dump cstatus_csv_dumper_1438;
    df_fifo_monitor fifo_monitor_1438;
    df_fifo_intf fifo_intf_1439(clock,reset);
    assign fifo_intf_1439.rd_en = AESL_inst_myproject.layer3_out_86_U.if_read & AESL_inst_myproject.layer3_out_86_U.if_empty_n;
    assign fifo_intf_1439.wr_en = AESL_inst_myproject.layer3_out_86_U.if_write & AESL_inst_myproject.layer3_out_86_U.if_full_n;
    assign fifo_intf_1439.fifo_rd_block = 0;
    assign fifo_intf_1439.fifo_wr_block = 0;
    assign fifo_intf_1439.finish = finish;
    csv_file_dump fifo_csv_dumper_1439;
    csv_file_dump cstatus_csv_dumper_1439;
    df_fifo_monitor fifo_monitor_1439;
    df_fifo_intf fifo_intf_1440(clock,reset);
    assign fifo_intf_1440.rd_en = AESL_inst_myproject.layer3_out_87_U.if_read & AESL_inst_myproject.layer3_out_87_U.if_empty_n;
    assign fifo_intf_1440.wr_en = AESL_inst_myproject.layer3_out_87_U.if_write & AESL_inst_myproject.layer3_out_87_U.if_full_n;
    assign fifo_intf_1440.fifo_rd_block = 0;
    assign fifo_intf_1440.fifo_wr_block = 0;
    assign fifo_intf_1440.finish = finish;
    csv_file_dump fifo_csv_dumper_1440;
    csv_file_dump cstatus_csv_dumper_1440;
    df_fifo_monitor fifo_monitor_1440;
    df_fifo_intf fifo_intf_1441(clock,reset);
    assign fifo_intf_1441.rd_en = AESL_inst_myproject.layer3_out_88_U.if_read & AESL_inst_myproject.layer3_out_88_U.if_empty_n;
    assign fifo_intf_1441.wr_en = AESL_inst_myproject.layer3_out_88_U.if_write & AESL_inst_myproject.layer3_out_88_U.if_full_n;
    assign fifo_intf_1441.fifo_rd_block = 0;
    assign fifo_intf_1441.fifo_wr_block = 0;
    assign fifo_intf_1441.finish = finish;
    csv_file_dump fifo_csv_dumper_1441;
    csv_file_dump cstatus_csv_dumper_1441;
    df_fifo_monitor fifo_monitor_1441;
    df_fifo_intf fifo_intf_1442(clock,reset);
    assign fifo_intf_1442.rd_en = AESL_inst_myproject.layer3_out_89_U.if_read & AESL_inst_myproject.layer3_out_89_U.if_empty_n;
    assign fifo_intf_1442.wr_en = AESL_inst_myproject.layer3_out_89_U.if_write & AESL_inst_myproject.layer3_out_89_U.if_full_n;
    assign fifo_intf_1442.fifo_rd_block = 0;
    assign fifo_intf_1442.fifo_wr_block = 0;
    assign fifo_intf_1442.finish = finish;
    csv_file_dump fifo_csv_dumper_1442;
    csv_file_dump cstatus_csv_dumper_1442;
    df_fifo_monitor fifo_monitor_1442;
    df_fifo_intf fifo_intf_1443(clock,reset);
    assign fifo_intf_1443.rd_en = AESL_inst_myproject.layer3_out_90_U.if_read & AESL_inst_myproject.layer3_out_90_U.if_empty_n;
    assign fifo_intf_1443.wr_en = AESL_inst_myproject.layer3_out_90_U.if_write & AESL_inst_myproject.layer3_out_90_U.if_full_n;
    assign fifo_intf_1443.fifo_rd_block = 0;
    assign fifo_intf_1443.fifo_wr_block = 0;
    assign fifo_intf_1443.finish = finish;
    csv_file_dump fifo_csv_dumper_1443;
    csv_file_dump cstatus_csv_dumper_1443;
    df_fifo_monitor fifo_monitor_1443;
    df_fifo_intf fifo_intf_1444(clock,reset);
    assign fifo_intf_1444.rd_en = AESL_inst_myproject.layer3_out_91_U.if_read & AESL_inst_myproject.layer3_out_91_U.if_empty_n;
    assign fifo_intf_1444.wr_en = AESL_inst_myproject.layer3_out_91_U.if_write & AESL_inst_myproject.layer3_out_91_U.if_full_n;
    assign fifo_intf_1444.fifo_rd_block = 0;
    assign fifo_intf_1444.fifo_wr_block = 0;
    assign fifo_intf_1444.finish = finish;
    csv_file_dump fifo_csv_dumper_1444;
    csv_file_dump cstatus_csv_dumper_1444;
    df_fifo_monitor fifo_monitor_1444;
    df_fifo_intf fifo_intf_1445(clock,reset);
    assign fifo_intf_1445.rd_en = AESL_inst_myproject.layer3_out_92_U.if_read & AESL_inst_myproject.layer3_out_92_U.if_empty_n;
    assign fifo_intf_1445.wr_en = AESL_inst_myproject.layer3_out_92_U.if_write & AESL_inst_myproject.layer3_out_92_U.if_full_n;
    assign fifo_intf_1445.fifo_rd_block = 0;
    assign fifo_intf_1445.fifo_wr_block = 0;
    assign fifo_intf_1445.finish = finish;
    csv_file_dump fifo_csv_dumper_1445;
    csv_file_dump cstatus_csv_dumper_1445;
    df_fifo_monitor fifo_monitor_1445;
    df_fifo_intf fifo_intf_1446(clock,reset);
    assign fifo_intf_1446.rd_en = AESL_inst_myproject.layer3_out_93_U.if_read & AESL_inst_myproject.layer3_out_93_U.if_empty_n;
    assign fifo_intf_1446.wr_en = AESL_inst_myproject.layer3_out_93_U.if_write & AESL_inst_myproject.layer3_out_93_U.if_full_n;
    assign fifo_intf_1446.fifo_rd_block = 0;
    assign fifo_intf_1446.fifo_wr_block = 0;
    assign fifo_intf_1446.finish = finish;
    csv_file_dump fifo_csv_dumper_1446;
    csv_file_dump cstatus_csv_dumper_1446;
    df_fifo_monitor fifo_monitor_1446;
    df_fifo_intf fifo_intf_1447(clock,reset);
    assign fifo_intf_1447.rd_en = AESL_inst_myproject.layer3_out_94_U.if_read & AESL_inst_myproject.layer3_out_94_U.if_empty_n;
    assign fifo_intf_1447.wr_en = AESL_inst_myproject.layer3_out_94_U.if_write & AESL_inst_myproject.layer3_out_94_U.if_full_n;
    assign fifo_intf_1447.fifo_rd_block = 0;
    assign fifo_intf_1447.fifo_wr_block = 0;
    assign fifo_intf_1447.finish = finish;
    csv_file_dump fifo_csv_dumper_1447;
    csv_file_dump cstatus_csv_dumper_1447;
    df_fifo_monitor fifo_monitor_1447;
    df_fifo_intf fifo_intf_1448(clock,reset);
    assign fifo_intf_1448.rd_en = AESL_inst_myproject.layer3_out_95_U.if_read & AESL_inst_myproject.layer3_out_95_U.if_empty_n;
    assign fifo_intf_1448.wr_en = AESL_inst_myproject.layer3_out_95_U.if_write & AESL_inst_myproject.layer3_out_95_U.if_full_n;
    assign fifo_intf_1448.fifo_rd_block = 0;
    assign fifo_intf_1448.fifo_wr_block = 0;
    assign fifo_intf_1448.finish = finish;
    csv_file_dump fifo_csv_dumper_1448;
    csv_file_dump cstatus_csv_dumper_1448;
    df_fifo_monitor fifo_monitor_1448;
    df_fifo_intf fifo_intf_1449(clock,reset);
    assign fifo_intf_1449.rd_en = AESL_inst_myproject.layer3_out_96_U.if_read & AESL_inst_myproject.layer3_out_96_U.if_empty_n;
    assign fifo_intf_1449.wr_en = AESL_inst_myproject.layer3_out_96_U.if_write & AESL_inst_myproject.layer3_out_96_U.if_full_n;
    assign fifo_intf_1449.fifo_rd_block = 0;
    assign fifo_intf_1449.fifo_wr_block = 0;
    assign fifo_intf_1449.finish = finish;
    csv_file_dump fifo_csv_dumper_1449;
    csv_file_dump cstatus_csv_dumper_1449;
    df_fifo_monitor fifo_monitor_1449;
    df_fifo_intf fifo_intf_1450(clock,reset);
    assign fifo_intf_1450.rd_en = AESL_inst_myproject.layer3_out_97_U.if_read & AESL_inst_myproject.layer3_out_97_U.if_empty_n;
    assign fifo_intf_1450.wr_en = AESL_inst_myproject.layer3_out_97_U.if_write & AESL_inst_myproject.layer3_out_97_U.if_full_n;
    assign fifo_intf_1450.fifo_rd_block = 0;
    assign fifo_intf_1450.fifo_wr_block = 0;
    assign fifo_intf_1450.finish = finish;
    csv_file_dump fifo_csv_dumper_1450;
    csv_file_dump cstatus_csv_dumper_1450;
    df_fifo_monitor fifo_monitor_1450;
    df_fifo_intf fifo_intf_1451(clock,reset);
    assign fifo_intf_1451.rd_en = AESL_inst_myproject.layer3_out_98_U.if_read & AESL_inst_myproject.layer3_out_98_U.if_empty_n;
    assign fifo_intf_1451.wr_en = AESL_inst_myproject.layer3_out_98_U.if_write & AESL_inst_myproject.layer3_out_98_U.if_full_n;
    assign fifo_intf_1451.fifo_rd_block = 0;
    assign fifo_intf_1451.fifo_wr_block = 0;
    assign fifo_intf_1451.finish = finish;
    csv_file_dump fifo_csv_dumper_1451;
    csv_file_dump cstatus_csv_dumper_1451;
    df_fifo_monitor fifo_monitor_1451;
    df_fifo_intf fifo_intf_1452(clock,reset);
    assign fifo_intf_1452.rd_en = AESL_inst_myproject.layer3_out_99_U.if_read & AESL_inst_myproject.layer3_out_99_U.if_empty_n;
    assign fifo_intf_1452.wr_en = AESL_inst_myproject.layer3_out_99_U.if_write & AESL_inst_myproject.layer3_out_99_U.if_full_n;
    assign fifo_intf_1452.fifo_rd_block = 0;
    assign fifo_intf_1452.fifo_wr_block = 0;
    assign fifo_intf_1452.finish = finish;
    csv_file_dump fifo_csv_dumper_1452;
    csv_file_dump cstatus_csv_dumper_1452;
    df_fifo_monitor fifo_monitor_1452;
    df_fifo_intf fifo_intf_1453(clock,reset);
    assign fifo_intf_1453.rd_en = AESL_inst_myproject.layer3_out_100_U.if_read & AESL_inst_myproject.layer3_out_100_U.if_empty_n;
    assign fifo_intf_1453.wr_en = AESL_inst_myproject.layer3_out_100_U.if_write & AESL_inst_myproject.layer3_out_100_U.if_full_n;
    assign fifo_intf_1453.fifo_rd_block = 0;
    assign fifo_intf_1453.fifo_wr_block = 0;
    assign fifo_intf_1453.finish = finish;
    csv_file_dump fifo_csv_dumper_1453;
    csv_file_dump cstatus_csv_dumper_1453;
    df_fifo_monitor fifo_monitor_1453;
    df_fifo_intf fifo_intf_1454(clock,reset);
    assign fifo_intf_1454.rd_en = AESL_inst_myproject.layer3_out_101_U.if_read & AESL_inst_myproject.layer3_out_101_U.if_empty_n;
    assign fifo_intf_1454.wr_en = AESL_inst_myproject.layer3_out_101_U.if_write & AESL_inst_myproject.layer3_out_101_U.if_full_n;
    assign fifo_intf_1454.fifo_rd_block = 0;
    assign fifo_intf_1454.fifo_wr_block = 0;
    assign fifo_intf_1454.finish = finish;
    csv_file_dump fifo_csv_dumper_1454;
    csv_file_dump cstatus_csv_dumper_1454;
    df_fifo_monitor fifo_monitor_1454;
    df_fifo_intf fifo_intf_1455(clock,reset);
    assign fifo_intf_1455.rd_en = AESL_inst_myproject.layer3_out_102_U.if_read & AESL_inst_myproject.layer3_out_102_U.if_empty_n;
    assign fifo_intf_1455.wr_en = AESL_inst_myproject.layer3_out_102_U.if_write & AESL_inst_myproject.layer3_out_102_U.if_full_n;
    assign fifo_intf_1455.fifo_rd_block = 0;
    assign fifo_intf_1455.fifo_wr_block = 0;
    assign fifo_intf_1455.finish = finish;
    csv_file_dump fifo_csv_dumper_1455;
    csv_file_dump cstatus_csv_dumper_1455;
    df_fifo_monitor fifo_monitor_1455;
    df_fifo_intf fifo_intf_1456(clock,reset);
    assign fifo_intf_1456.rd_en = AESL_inst_myproject.layer3_out_103_U.if_read & AESL_inst_myproject.layer3_out_103_U.if_empty_n;
    assign fifo_intf_1456.wr_en = AESL_inst_myproject.layer3_out_103_U.if_write & AESL_inst_myproject.layer3_out_103_U.if_full_n;
    assign fifo_intf_1456.fifo_rd_block = 0;
    assign fifo_intf_1456.fifo_wr_block = 0;
    assign fifo_intf_1456.finish = finish;
    csv_file_dump fifo_csv_dumper_1456;
    csv_file_dump cstatus_csv_dumper_1456;
    df_fifo_monitor fifo_monitor_1456;
    df_fifo_intf fifo_intf_1457(clock,reset);
    assign fifo_intf_1457.rd_en = AESL_inst_myproject.layer3_out_104_U.if_read & AESL_inst_myproject.layer3_out_104_U.if_empty_n;
    assign fifo_intf_1457.wr_en = AESL_inst_myproject.layer3_out_104_U.if_write & AESL_inst_myproject.layer3_out_104_U.if_full_n;
    assign fifo_intf_1457.fifo_rd_block = 0;
    assign fifo_intf_1457.fifo_wr_block = 0;
    assign fifo_intf_1457.finish = finish;
    csv_file_dump fifo_csv_dumper_1457;
    csv_file_dump cstatus_csv_dumper_1457;
    df_fifo_monitor fifo_monitor_1457;
    df_fifo_intf fifo_intf_1458(clock,reset);
    assign fifo_intf_1458.rd_en = AESL_inst_myproject.layer3_out_105_U.if_read & AESL_inst_myproject.layer3_out_105_U.if_empty_n;
    assign fifo_intf_1458.wr_en = AESL_inst_myproject.layer3_out_105_U.if_write & AESL_inst_myproject.layer3_out_105_U.if_full_n;
    assign fifo_intf_1458.fifo_rd_block = 0;
    assign fifo_intf_1458.fifo_wr_block = 0;
    assign fifo_intf_1458.finish = finish;
    csv_file_dump fifo_csv_dumper_1458;
    csv_file_dump cstatus_csv_dumper_1458;
    df_fifo_monitor fifo_monitor_1458;
    df_fifo_intf fifo_intf_1459(clock,reset);
    assign fifo_intf_1459.rd_en = AESL_inst_myproject.layer3_out_106_U.if_read & AESL_inst_myproject.layer3_out_106_U.if_empty_n;
    assign fifo_intf_1459.wr_en = AESL_inst_myproject.layer3_out_106_U.if_write & AESL_inst_myproject.layer3_out_106_U.if_full_n;
    assign fifo_intf_1459.fifo_rd_block = 0;
    assign fifo_intf_1459.fifo_wr_block = 0;
    assign fifo_intf_1459.finish = finish;
    csv_file_dump fifo_csv_dumper_1459;
    csv_file_dump cstatus_csv_dumper_1459;
    df_fifo_monitor fifo_monitor_1459;
    df_fifo_intf fifo_intf_1460(clock,reset);
    assign fifo_intf_1460.rd_en = AESL_inst_myproject.layer3_out_107_U.if_read & AESL_inst_myproject.layer3_out_107_U.if_empty_n;
    assign fifo_intf_1460.wr_en = AESL_inst_myproject.layer3_out_107_U.if_write & AESL_inst_myproject.layer3_out_107_U.if_full_n;
    assign fifo_intf_1460.fifo_rd_block = 0;
    assign fifo_intf_1460.fifo_wr_block = 0;
    assign fifo_intf_1460.finish = finish;
    csv_file_dump fifo_csv_dumper_1460;
    csv_file_dump cstatus_csv_dumper_1460;
    df_fifo_monitor fifo_monitor_1460;
    df_fifo_intf fifo_intf_1461(clock,reset);
    assign fifo_intf_1461.rd_en = AESL_inst_myproject.layer3_out_108_U.if_read & AESL_inst_myproject.layer3_out_108_U.if_empty_n;
    assign fifo_intf_1461.wr_en = AESL_inst_myproject.layer3_out_108_U.if_write & AESL_inst_myproject.layer3_out_108_U.if_full_n;
    assign fifo_intf_1461.fifo_rd_block = 0;
    assign fifo_intf_1461.fifo_wr_block = 0;
    assign fifo_intf_1461.finish = finish;
    csv_file_dump fifo_csv_dumper_1461;
    csv_file_dump cstatus_csv_dumper_1461;
    df_fifo_monitor fifo_monitor_1461;
    df_fifo_intf fifo_intf_1462(clock,reset);
    assign fifo_intf_1462.rd_en = AESL_inst_myproject.layer3_out_109_U.if_read & AESL_inst_myproject.layer3_out_109_U.if_empty_n;
    assign fifo_intf_1462.wr_en = AESL_inst_myproject.layer3_out_109_U.if_write & AESL_inst_myproject.layer3_out_109_U.if_full_n;
    assign fifo_intf_1462.fifo_rd_block = 0;
    assign fifo_intf_1462.fifo_wr_block = 0;
    assign fifo_intf_1462.finish = finish;
    csv_file_dump fifo_csv_dumper_1462;
    csv_file_dump cstatus_csv_dumper_1462;
    df_fifo_monitor fifo_monitor_1462;
    df_fifo_intf fifo_intf_1463(clock,reset);
    assign fifo_intf_1463.rd_en = AESL_inst_myproject.layer3_out_110_U.if_read & AESL_inst_myproject.layer3_out_110_U.if_empty_n;
    assign fifo_intf_1463.wr_en = AESL_inst_myproject.layer3_out_110_U.if_write & AESL_inst_myproject.layer3_out_110_U.if_full_n;
    assign fifo_intf_1463.fifo_rd_block = 0;
    assign fifo_intf_1463.fifo_wr_block = 0;
    assign fifo_intf_1463.finish = finish;
    csv_file_dump fifo_csv_dumper_1463;
    csv_file_dump cstatus_csv_dumper_1463;
    df_fifo_monitor fifo_monitor_1463;
    df_fifo_intf fifo_intf_1464(clock,reset);
    assign fifo_intf_1464.rd_en = AESL_inst_myproject.layer3_out_111_U.if_read & AESL_inst_myproject.layer3_out_111_U.if_empty_n;
    assign fifo_intf_1464.wr_en = AESL_inst_myproject.layer3_out_111_U.if_write & AESL_inst_myproject.layer3_out_111_U.if_full_n;
    assign fifo_intf_1464.fifo_rd_block = 0;
    assign fifo_intf_1464.fifo_wr_block = 0;
    assign fifo_intf_1464.finish = finish;
    csv_file_dump fifo_csv_dumper_1464;
    csv_file_dump cstatus_csv_dumper_1464;
    df_fifo_monitor fifo_monitor_1464;
    df_fifo_intf fifo_intf_1465(clock,reset);
    assign fifo_intf_1465.rd_en = AESL_inst_myproject.layer3_out_112_U.if_read & AESL_inst_myproject.layer3_out_112_U.if_empty_n;
    assign fifo_intf_1465.wr_en = AESL_inst_myproject.layer3_out_112_U.if_write & AESL_inst_myproject.layer3_out_112_U.if_full_n;
    assign fifo_intf_1465.fifo_rd_block = 0;
    assign fifo_intf_1465.fifo_wr_block = 0;
    assign fifo_intf_1465.finish = finish;
    csv_file_dump fifo_csv_dumper_1465;
    csv_file_dump cstatus_csv_dumper_1465;
    df_fifo_monitor fifo_monitor_1465;
    df_fifo_intf fifo_intf_1466(clock,reset);
    assign fifo_intf_1466.rd_en = AESL_inst_myproject.layer3_out_113_U.if_read & AESL_inst_myproject.layer3_out_113_U.if_empty_n;
    assign fifo_intf_1466.wr_en = AESL_inst_myproject.layer3_out_113_U.if_write & AESL_inst_myproject.layer3_out_113_U.if_full_n;
    assign fifo_intf_1466.fifo_rd_block = 0;
    assign fifo_intf_1466.fifo_wr_block = 0;
    assign fifo_intf_1466.finish = finish;
    csv_file_dump fifo_csv_dumper_1466;
    csv_file_dump cstatus_csv_dumper_1466;
    df_fifo_monitor fifo_monitor_1466;
    df_fifo_intf fifo_intf_1467(clock,reset);
    assign fifo_intf_1467.rd_en = AESL_inst_myproject.layer3_out_114_U.if_read & AESL_inst_myproject.layer3_out_114_U.if_empty_n;
    assign fifo_intf_1467.wr_en = AESL_inst_myproject.layer3_out_114_U.if_write & AESL_inst_myproject.layer3_out_114_U.if_full_n;
    assign fifo_intf_1467.fifo_rd_block = 0;
    assign fifo_intf_1467.fifo_wr_block = 0;
    assign fifo_intf_1467.finish = finish;
    csv_file_dump fifo_csv_dumper_1467;
    csv_file_dump cstatus_csv_dumper_1467;
    df_fifo_monitor fifo_monitor_1467;
    df_fifo_intf fifo_intf_1468(clock,reset);
    assign fifo_intf_1468.rd_en = AESL_inst_myproject.layer3_out_115_U.if_read & AESL_inst_myproject.layer3_out_115_U.if_empty_n;
    assign fifo_intf_1468.wr_en = AESL_inst_myproject.layer3_out_115_U.if_write & AESL_inst_myproject.layer3_out_115_U.if_full_n;
    assign fifo_intf_1468.fifo_rd_block = 0;
    assign fifo_intf_1468.fifo_wr_block = 0;
    assign fifo_intf_1468.finish = finish;
    csv_file_dump fifo_csv_dumper_1468;
    csv_file_dump cstatus_csv_dumper_1468;
    df_fifo_monitor fifo_monitor_1468;
    df_fifo_intf fifo_intf_1469(clock,reset);
    assign fifo_intf_1469.rd_en = AESL_inst_myproject.layer3_out_116_U.if_read & AESL_inst_myproject.layer3_out_116_U.if_empty_n;
    assign fifo_intf_1469.wr_en = AESL_inst_myproject.layer3_out_116_U.if_write & AESL_inst_myproject.layer3_out_116_U.if_full_n;
    assign fifo_intf_1469.fifo_rd_block = 0;
    assign fifo_intf_1469.fifo_wr_block = 0;
    assign fifo_intf_1469.finish = finish;
    csv_file_dump fifo_csv_dumper_1469;
    csv_file_dump cstatus_csv_dumper_1469;
    df_fifo_monitor fifo_monitor_1469;
    df_fifo_intf fifo_intf_1470(clock,reset);
    assign fifo_intf_1470.rd_en = AESL_inst_myproject.layer3_out_117_U.if_read & AESL_inst_myproject.layer3_out_117_U.if_empty_n;
    assign fifo_intf_1470.wr_en = AESL_inst_myproject.layer3_out_117_U.if_write & AESL_inst_myproject.layer3_out_117_U.if_full_n;
    assign fifo_intf_1470.fifo_rd_block = 0;
    assign fifo_intf_1470.fifo_wr_block = 0;
    assign fifo_intf_1470.finish = finish;
    csv_file_dump fifo_csv_dumper_1470;
    csv_file_dump cstatus_csv_dumper_1470;
    df_fifo_monitor fifo_monitor_1470;
    df_fifo_intf fifo_intf_1471(clock,reset);
    assign fifo_intf_1471.rd_en = AESL_inst_myproject.layer3_out_118_U.if_read & AESL_inst_myproject.layer3_out_118_U.if_empty_n;
    assign fifo_intf_1471.wr_en = AESL_inst_myproject.layer3_out_118_U.if_write & AESL_inst_myproject.layer3_out_118_U.if_full_n;
    assign fifo_intf_1471.fifo_rd_block = 0;
    assign fifo_intf_1471.fifo_wr_block = 0;
    assign fifo_intf_1471.finish = finish;
    csv_file_dump fifo_csv_dumper_1471;
    csv_file_dump cstatus_csv_dumper_1471;
    df_fifo_monitor fifo_monitor_1471;
    df_fifo_intf fifo_intf_1472(clock,reset);
    assign fifo_intf_1472.rd_en = AESL_inst_myproject.layer3_out_119_U.if_read & AESL_inst_myproject.layer3_out_119_U.if_empty_n;
    assign fifo_intf_1472.wr_en = AESL_inst_myproject.layer3_out_119_U.if_write & AESL_inst_myproject.layer3_out_119_U.if_full_n;
    assign fifo_intf_1472.fifo_rd_block = 0;
    assign fifo_intf_1472.fifo_wr_block = 0;
    assign fifo_intf_1472.finish = finish;
    csv_file_dump fifo_csv_dumper_1472;
    csv_file_dump cstatus_csv_dumper_1472;
    df_fifo_monitor fifo_monitor_1472;
    df_fifo_intf fifo_intf_1473(clock,reset);
    assign fifo_intf_1473.rd_en = AESL_inst_myproject.layer3_out_120_U.if_read & AESL_inst_myproject.layer3_out_120_U.if_empty_n;
    assign fifo_intf_1473.wr_en = AESL_inst_myproject.layer3_out_120_U.if_write & AESL_inst_myproject.layer3_out_120_U.if_full_n;
    assign fifo_intf_1473.fifo_rd_block = 0;
    assign fifo_intf_1473.fifo_wr_block = 0;
    assign fifo_intf_1473.finish = finish;
    csv_file_dump fifo_csv_dumper_1473;
    csv_file_dump cstatus_csv_dumper_1473;
    df_fifo_monitor fifo_monitor_1473;
    df_fifo_intf fifo_intf_1474(clock,reset);
    assign fifo_intf_1474.rd_en = AESL_inst_myproject.layer3_out_121_U.if_read & AESL_inst_myproject.layer3_out_121_U.if_empty_n;
    assign fifo_intf_1474.wr_en = AESL_inst_myproject.layer3_out_121_U.if_write & AESL_inst_myproject.layer3_out_121_U.if_full_n;
    assign fifo_intf_1474.fifo_rd_block = 0;
    assign fifo_intf_1474.fifo_wr_block = 0;
    assign fifo_intf_1474.finish = finish;
    csv_file_dump fifo_csv_dumper_1474;
    csv_file_dump cstatus_csv_dumper_1474;
    df_fifo_monitor fifo_monitor_1474;
    df_fifo_intf fifo_intf_1475(clock,reset);
    assign fifo_intf_1475.rd_en = AESL_inst_myproject.layer3_out_122_U.if_read & AESL_inst_myproject.layer3_out_122_U.if_empty_n;
    assign fifo_intf_1475.wr_en = AESL_inst_myproject.layer3_out_122_U.if_write & AESL_inst_myproject.layer3_out_122_U.if_full_n;
    assign fifo_intf_1475.fifo_rd_block = 0;
    assign fifo_intf_1475.fifo_wr_block = 0;
    assign fifo_intf_1475.finish = finish;
    csv_file_dump fifo_csv_dumper_1475;
    csv_file_dump cstatus_csv_dumper_1475;
    df_fifo_monitor fifo_monitor_1475;
    df_fifo_intf fifo_intf_1476(clock,reset);
    assign fifo_intf_1476.rd_en = AESL_inst_myproject.layer3_out_123_U.if_read & AESL_inst_myproject.layer3_out_123_U.if_empty_n;
    assign fifo_intf_1476.wr_en = AESL_inst_myproject.layer3_out_123_U.if_write & AESL_inst_myproject.layer3_out_123_U.if_full_n;
    assign fifo_intf_1476.fifo_rd_block = 0;
    assign fifo_intf_1476.fifo_wr_block = 0;
    assign fifo_intf_1476.finish = finish;
    csv_file_dump fifo_csv_dumper_1476;
    csv_file_dump cstatus_csv_dumper_1476;
    df_fifo_monitor fifo_monitor_1476;
    df_fifo_intf fifo_intf_1477(clock,reset);
    assign fifo_intf_1477.rd_en = AESL_inst_myproject.layer3_out_124_U.if_read & AESL_inst_myproject.layer3_out_124_U.if_empty_n;
    assign fifo_intf_1477.wr_en = AESL_inst_myproject.layer3_out_124_U.if_write & AESL_inst_myproject.layer3_out_124_U.if_full_n;
    assign fifo_intf_1477.fifo_rd_block = 0;
    assign fifo_intf_1477.fifo_wr_block = 0;
    assign fifo_intf_1477.finish = finish;
    csv_file_dump fifo_csv_dumper_1477;
    csv_file_dump cstatus_csv_dumper_1477;
    df_fifo_monitor fifo_monitor_1477;
    df_fifo_intf fifo_intf_1478(clock,reset);
    assign fifo_intf_1478.rd_en = AESL_inst_myproject.layer3_out_125_U.if_read & AESL_inst_myproject.layer3_out_125_U.if_empty_n;
    assign fifo_intf_1478.wr_en = AESL_inst_myproject.layer3_out_125_U.if_write & AESL_inst_myproject.layer3_out_125_U.if_full_n;
    assign fifo_intf_1478.fifo_rd_block = 0;
    assign fifo_intf_1478.fifo_wr_block = 0;
    assign fifo_intf_1478.finish = finish;
    csv_file_dump fifo_csv_dumper_1478;
    csv_file_dump cstatus_csv_dumper_1478;
    df_fifo_monitor fifo_monitor_1478;
    df_fifo_intf fifo_intf_1479(clock,reset);
    assign fifo_intf_1479.rd_en = AESL_inst_myproject.layer3_out_126_U.if_read & AESL_inst_myproject.layer3_out_126_U.if_empty_n;
    assign fifo_intf_1479.wr_en = AESL_inst_myproject.layer3_out_126_U.if_write & AESL_inst_myproject.layer3_out_126_U.if_full_n;
    assign fifo_intf_1479.fifo_rd_block = 0;
    assign fifo_intf_1479.fifo_wr_block = 0;
    assign fifo_intf_1479.finish = finish;
    csv_file_dump fifo_csv_dumper_1479;
    csv_file_dump cstatus_csv_dumper_1479;
    df_fifo_monitor fifo_monitor_1479;
    df_fifo_intf fifo_intf_1480(clock,reset);
    assign fifo_intf_1480.rd_en = AESL_inst_myproject.layer3_out_127_U.if_read & AESL_inst_myproject.layer3_out_127_U.if_empty_n;
    assign fifo_intf_1480.wr_en = AESL_inst_myproject.layer3_out_127_U.if_write & AESL_inst_myproject.layer3_out_127_U.if_full_n;
    assign fifo_intf_1480.fifo_rd_block = 0;
    assign fifo_intf_1480.fifo_wr_block = 0;
    assign fifo_intf_1480.finish = finish;
    csv_file_dump fifo_csv_dumper_1480;
    csv_file_dump cstatus_csv_dumper_1480;
    df_fifo_monitor fifo_monitor_1480;
    df_fifo_intf fifo_intf_1481(clock,reset);
    assign fifo_intf_1481.rd_en = AESL_inst_myproject.layer3_out_128_U.if_read & AESL_inst_myproject.layer3_out_128_U.if_empty_n;
    assign fifo_intf_1481.wr_en = AESL_inst_myproject.layer3_out_128_U.if_write & AESL_inst_myproject.layer3_out_128_U.if_full_n;
    assign fifo_intf_1481.fifo_rd_block = 0;
    assign fifo_intf_1481.fifo_wr_block = 0;
    assign fifo_intf_1481.finish = finish;
    csv_file_dump fifo_csv_dumper_1481;
    csv_file_dump cstatus_csv_dumper_1481;
    df_fifo_monitor fifo_monitor_1481;
    df_fifo_intf fifo_intf_1482(clock,reset);
    assign fifo_intf_1482.rd_en = AESL_inst_myproject.layer3_out_129_U.if_read & AESL_inst_myproject.layer3_out_129_U.if_empty_n;
    assign fifo_intf_1482.wr_en = AESL_inst_myproject.layer3_out_129_U.if_write & AESL_inst_myproject.layer3_out_129_U.if_full_n;
    assign fifo_intf_1482.fifo_rd_block = 0;
    assign fifo_intf_1482.fifo_wr_block = 0;
    assign fifo_intf_1482.finish = finish;
    csv_file_dump fifo_csv_dumper_1482;
    csv_file_dump cstatus_csv_dumper_1482;
    df_fifo_monitor fifo_monitor_1482;
    df_fifo_intf fifo_intf_1483(clock,reset);
    assign fifo_intf_1483.rd_en = AESL_inst_myproject.layer3_out_130_U.if_read & AESL_inst_myproject.layer3_out_130_U.if_empty_n;
    assign fifo_intf_1483.wr_en = AESL_inst_myproject.layer3_out_130_U.if_write & AESL_inst_myproject.layer3_out_130_U.if_full_n;
    assign fifo_intf_1483.fifo_rd_block = 0;
    assign fifo_intf_1483.fifo_wr_block = 0;
    assign fifo_intf_1483.finish = finish;
    csv_file_dump fifo_csv_dumper_1483;
    csv_file_dump cstatus_csv_dumper_1483;
    df_fifo_monitor fifo_monitor_1483;
    df_fifo_intf fifo_intf_1484(clock,reset);
    assign fifo_intf_1484.rd_en = AESL_inst_myproject.layer3_out_131_U.if_read & AESL_inst_myproject.layer3_out_131_U.if_empty_n;
    assign fifo_intf_1484.wr_en = AESL_inst_myproject.layer3_out_131_U.if_write & AESL_inst_myproject.layer3_out_131_U.if_full_n;
    assign fifo_intf_1484.fifo_rd_block = 0;
    assign fifo_intf_1484.fifo_wr_block = 0;
    assign fifo_intf_1484.finish = finish;
    csv_file_dump fifo_csv_dumper_1484;
    csv_file_dump cstatus_csv_dumper_1484;
    df_fifo_monitor fifo_monitor_1484;
    df_fifo_intf fifo_intf_1485(clock,reset);
    assign fifo_intf_1485.rd_en = AESL_inst_myproject.layer3_out_132_U.if_read & AESL_inst_myproject.layer3_out_132_U.if_empty_n;
    assign fifo_intf_1485.wr_en = AESL_inst_myproject.layer3_out_132_U.if_write & AESL_inst_myproject.layer3_out_132_U.if_full_n;
    assign fifo_intf_1485.fifo_rd_block = 0;
    assign fifo_intf_1485.fifo_wr_block = 0;
    assign fifo_intf_1485.finish = finish;
    csv_file_dump fifo_csv_dumper_1485;
    csv_file_dump cstatus_csv_dumper_1485;
    df_fifo_monitor fifo_monitor_1485;
    df_fifo_intf fifo_intf_1486(clock,reset);
    assign fifo_intf_1486.rd_en = AESL_inst_myproject.layer3_out_133_U.if_read & AESL_inst_myproject.layer3_out_133_U.if_empty_n;
    assign fifo_intf_1486.wr_en = AESL_inst_myproject.layer3_out_133_U.if_write & AESL_inst_myproject.layer3_out_133_U.if_full_n;
    assign fifo_intf_1486.fifo_rd_block = 0;
    assign fifo_intf_1486.fifo_wr_block = 0;
    assign fifo_intf_1486.finish = finish;
    csv_file_dump fifo_csv_dumper_1486;
    csv_file_dump cstatus_csv_dumper_1486;
    df_fifo_monitor fifo_monitor_1486;
    df_fifo_intf fifo_intf_1487(clock,reset);
    assign fifo_intf_1487.rd_en = AESL_inst_myproject.layer3_out_134_U.if_read & AESL_inst_myproject.layer3_out_134_U.if_empty_n;
    assign fifo_intf_1487.wr_en = AESL_inst_myproject.layer3_out_134_U.if_write & AESL_inst_myproject.layer3_out_134_U.if_full_n;
    assign fifo_intf_1487.fifo_rd_block = 0;
    assign fifo_intf_1487.fifo_wr_block = 0;
    assign fifo_intf_1487.finish = finish;
    csv_file_dump fifo_csv_dumper_1487;
    csv_file_dump cstatus_csv_dumper_1487;
    df_fifo_monitor fifo_monitor_1487;
    df_fifo_intf fifo_intf_1488(clock,reset);
    assign fifo_intf_1488.rd_en = AESL_inst_myproject.layer3_out_135_U.if_read & AESL_inst_myproject.layer3_out_135_U.if_empty_n;
    assign fifo_intf_1488.wr_en = AESL_inst_myproject.layer3_out_135_U.if_write & AESL_inst_myproject.layer3_out_135_U.if_full_n;
    assign fifo_intf_1488.fifo_rd_block = 0;
    assign fifo_intf_1488.fifo_wr_block = 0;
    assign fifo_intf_1488.finish = finish;
    csv_file_dump fifo_csv_dumper_1488;
    csv_file_dump cstatus_csv_dumper_1488;
    df_fifo_monitor fifo_monitor_1488;
    df_fifo_intf fifo_intf_1489(clock,reset);
    assign fifo_intf_1489.rd_en = AESL_inst_myproject.layer3_out_136_U.if_read & AESL_inst_myproject.layer3_out_136_U.if_empty_n;
    assign fifo_intf_1489.wr_en = AESL_inst_myproject.layer3_out_136_U.if_write & AESL_inst_myproject.layer3_out_136_U.if_full_n;
    assign fifo_intf_1489.fifo_rd_block = 0;
    assign fifo_intf_1489.fifo_wr_block = 0;
    assign fifo_intf_1489.finish = finish;
    csv_file_dump fifo_csv_dumper_1489;
    csv_file_dump cstatus_csv_dumper_1489;
    df_fifo_monitor fifo_monitor_1489;
    df_fifo_intf fifo_intf_1490(clock,reset);
    assign fifo_intf_1490.rd_en = AESL_inst_myproject.layer3_out_137_U.if_read & AESL_inst_myproject.layer3_out_137_U.if_empty_n;
    assign fifo_intf_1490.wr_en = AESL_inst_myproject.layer3_out_137_U.if_write & AESL_inst_myproject.layer3_out_137_U.if_full_n;
    assign fifo_intf_1490.fifo_rd_block = 0;
    assign fifo_intf_1490.fifo_wr_block = 0;
    assign fifo_intf_1490.finish = finish;
    csv_file_dump fifo_csv_dumper_1490;
    csv_file_dump cstatus_csv_dumper_1490;
    df_fifo_monitor fifo_monitor_1490;
    df_fifo_intf fifo_intf_1491(clock,reset);
    assign fifo_intf_1491.rd_en = AESL_inst_myproject.layer3_out_138_U.if_read & AESL_inst_myproject.layer3_out_138_U.if_empty_n;
    assign fifo_intf_1491.wr_en = AESL_inst_myproject.layer3_out_138_U.if_write & AESL_inst_myproject.layer3_out_138_U.if_full_n;
    assign fifo_intf_1491.fifo_rd_block = 0;
    assign fifo_intf_1491.fifo_wr_block = 0;
    assign fifo_intf_1491.finish = finish;
    csv_file_dump fifo_csv_dumper_1491;
    csv_file_dump cstatus_csv_dumper_1491;
    df_fifo_monitor fifo_monitor_1491;
    df_fifo_intf fifo_intf_1492(clock,reset);
    assign fifo_intf_1492.rd_en = AESL_inst_myproject.layer3_out_139_U.if_read & AESL_inst_myproject.layer3_out_139_U.if_empty_n;
    assign fifo_intf_1492.wr_en = AESL_inst_myproject.layer3_out_139_U.if_write & AESL_inst_myproject.layer3_out_139_U.if_full_n;
    assign fifo_intf_1492.fifo_rd_block = 0;
    assign fifo_intf_1492.fifo_wr_block = 0;
    assign fifo_intf_1492.finish = finish;
    csv_file_dump fifo_csv_dumper_1492;
    csv_file_dump cstatus_csv_dumper_1492;
    df_fifo_monitor fifo_monitor_1492;
    df_fifo_intf fifo_intf_1493(clock,reset);
    assign fifo_intf_1493.rd_en = AESL_inst_myproject.layer3_out_140_U.if_read & AESL_inst_myproject.layer3_out_140_U.if_empty_n;
    assign fifo_intf_1493.wr_en = AESL_inst_myproject.layer3_out_140_U.if_write & AESL_inst_myproject.layer3_out_140_U.if_full_n;
    assign fifo_intf_1493.fifo_rd_block = 0;
    assign fifo_intf_1493.fifo_wr_block = 0;
    assign fifo_intf_1493.finish = finish;
    csv_file_dump fifo_csv_dumper_1493;
    csv_file_dump cstatus_csv_dumper_1493;
    df_fifo_monitor fifo_monitor_1493;
    df_fifo_intf fifo_intf_1494(clock,reset);
    assign fifo_intf_1494.rd_en = AESL_inst_myproject.layer3_out_141_U.if_read & AESL_inst_myproject.layer3_out_141_U.if_empty_n;
    assign fifo_intf_1494.wr_en = AESL_inst_myproject.layer3_out_141_U.if_write & AESL_inst_myproject.layer3_out_141_U.if_full_n;
    assign fifo_intf_1494.fifo_rd_block = 0;
    assign fifo_intf_1494.fifo_wr_block = 0;
    assign fifo_intf_1494.finish = finish;
    csv_file_dump fifo_csv_dumper_1494;
    csv_file_dump cstatus_csv_dumper_1494;
    df_fifo_monitor fifo_monitor_1494;
    df_fifo_intf fifo_intf_1495(clock,reset);
    assign fifo_intf_1495.rd_en = AESL_inst_myproject.layer3_out_142_U.if_read & AESL_inst_myproject.layer3_out_142_U.if_empty_n;
    assign fifo_intf_1495.wr_en = AESL_inst_myproject.layer3_out_142_U.if_write & AESL_inst_myproject.layer3_out_142_U.if_full_n;
    assign fifo_intf_1495.fifo_rd_block = 0;
    assign fifo_intf_1495.fifo_wr_block = 0;
    assign fifo_intf_1495.finish = finish;
    csv_file_dump fifo_csv_dumper_1495;
    csv_file_dump cstatus_csv_dumper_1495;
    df_fifo_monitor fifo_monitor_1495;
    df_fifo_intf fifo_intf_1496(clock,reset);
    assign fifo_intf_1496.rd_en = AESL_inst_myproject.layer3_out_143_U.if_read & AESL_inst_myproject.layer3_out_143_U.if_empty_n;
    assign fifo_intf_1496.wr_en = AESL_inst_myproject.layer3_out_143_U.if_write & AESL_inst_myproject.layer3_out_143_U.if_full_n;
    assign fifo_intf_1496.fifo_rd_block = 0;
    assign fifo_intf_1496.fifo_wr_block = 0;
    assign fifo_intf_1496.finish = finish;
    csv_file_dump fifo_csv_dumper_1496;
    csv_file_dump cstatus_csv_dumper_1496;
    df_fifo_monitor fifo_monitor_1496;
    df_fifo_intf fifo_intf_1497(clock,reset);
    assign fifo_intf_1497.rd_en = AESL_inst_myproject.layer3_out_144_U.if_read & AESL_inst_myproject.layer3_out_144_U.if_empty_n;
    assign fifo_intf_1497.wr_en = AESL_inst_myproject.layer3_out_144_U.if_write & AESL_inst_myproject.layer3_out_144_U.if_full_n;
    assign fifo_intf_1497.fifo_rd_block = 0;
    assign fifo_intf_1497.fifo_wr_block = 0;
    assign fifo_intf_1497.finish = finish;
    csv_file_dump fifo_csv_dumper_1497;
    csv_file_dump cstatus_csv_dumper_1497;
    df_fifo_monitor fifo_monitor_1497;
    df_fifo_intf fifo_intf_1498(clock,reset);
    assign fifo_intf_1498.rd_en = AESL_inst_myproject.layer3_out_145_U.if_read & AESL_inst_myproject.layer3_out_145_U.if_empty_n;
    assign fifo_intf_1498.wr_en = AESL_inst_myproject.layer3_out_145_U.if_write & AESL_inst_myproject.layer3_out_145_U.if_full_n;
    assign fifo_intf_1498.fifo_rd_block = 0;
    assign fifo_intf_1498.fifo_wr_block = 0;
    assign fifo_intf_1498.finish = finish;
    csv_file_dump fifo_csv_dumper_1498;
    csv_file_dump cstatus_csv_dumper_1498;
    df_fifo_monitor fifo_monitor_1498;
    df_fifo_intf fifo_intf_1499(clock,reset);
    assign fifo_intf_1499.rd_en = AESL_inst_myproject.layer3_out_146_U.if_read & AESL_inst_myproject.layer3_out_146_U.if_empty_n;
    assign fifo_intf_1499.wr_en = AESL_inst_myproject.layer3_out_146_U.if_write & AESL_inst_myproject.layer3_out_146_U.if_full_n;
    assign fifo_intf_1499.fifo_rd_block = 0;
    assign fifo_intf_1499.fifo_wr_block = 0;
    assign fifo_intf_1499.finish = finish;
    csv_file_dump fifo_csv_dumper_1499;
    csv_file_dump cstatus_csv_dumper_1499;
    df_fifo_monitor fifo_monitor_1499;
    df_fifo_intf fifo_intf_1500(clock,reset);
    assign fifo_intf_1500.rd_en = AESL_inst_myproject.layer3_out_147_U.if_read & AESL_inst_myproject.layer3_out_147_U.if_empty_n;
    assign fifo_intf_1500.wr_en = AESL_inst_myproject.layer3_out_147_U.if_write & AESL_inst_myproject.layer3_out_147_U.if_full_n;
    assign fifo_intf_1500.fifo_rd_block = 0;
    assign fifo_intf_1500.fifo_wr_block = 0;
    assign fifo_intf_1500.finish = finish;
    csv_file_dump fifo_csv_dumper_1500;
    csv_file_dump cstatus_csv_dumper_1500;
    df_fifo_monitor fifo_monitor_1500;
    df_fifo_intf fifo_intf_1501(clock,reset);
    assign fifo_intf_1501.rd_en = AESL_inst_myproject.layer3_out_148_U.if_read & AESL_inst_myproject.layer3_out_148_U.if_empty_n;
    assign fifo_intf_1501.wr_en = AESL_inst_myproject.layer3_out_148_U.if_write & AESL_inst_myproject.layer3_out_148_U.if_full_n;
    assign fifo_intf_1501.fifo_rd_block = 0;
    assign fifo_intf_1501.fifo_wr_block = 0;
    assign fifo_intf_1501.finish = finish;
    csv_file_dump fifo_csv_dumper_1501;
    csv_file_dump cstatus_csv_dumper_1501;
    df_fifo_monitor fifo_monitor_1501;
    df_fifo_intf fifo_intf_1502(clock,reset);
    assign fifo_intf_1502.rd_en = AESL_inst_myproject.layer3_out_149_U.if_read & AESL_inst_myproject.layer3_out_149_U.if_empty_n;
    assign fifo_intf_1502.wr_en = AESL_inst_myproject.layer3_out_149_U.if_write & AESL_inst_myproject.layer3_out_149_U.if_full_n;
    assign fifo_intf_1502.fifo_rd_block = 0;
    assign fifo_intf_1502.fifo_wr_block = 0;
    assign fifo_intf_1502.finish = finish;
    csv_file_dump fifo_csv_dumper_1502;
    csv_file_dump cstatus_csv_dumper_1502;
    df_fifo_monitor fifo_monitor_1502;
    df_fifo_intf fifo_intf_1503(clock,reset);
    assign fifo_intf_1503.rd_en = AESL_inst_myproject.layer3_out_150_U.if_read & AESL_inst_myproject.layer3_out_150_U.if_empty_n;
    assign fifo_intf_1503.wr_en = AESL_inst_myproject.layer3_out_150_U.if_write & AESL_inst_myproject.layer3_out_150_U.if_full_n;
    assign fifo_intf_1503.fifo_rd_block = 0;
    assign fifo_intf_1503.fifo_wr_block = 0;
    assign fifo_intf_1503.finish = finish;
    csv_file_dump fifo_csv_dumper_1503;
    csv_file_dump cstatus_csv_dumper_1503;
    df_fifo_monitor fifo_monitor_1503;
    df_fifo_intf fifo_intf_1504(clock,reset);
    assign fifo_intf_1504.rd_en = AESL_inst_myproject.layer3_out_151_U.if_read & AESL_inst_myproject.layer3_out_151_U.if_empty_n;
    assign fifo_intf_1504.wr_en = AESL_inst_myproject.layer3_out_151_U.if_write & AESL_inst_myproject.layer3_out_151_U.if_full_n;
    assign fifo_intf_1504.fifo_rd_block = 0;
    assign fifo_intf_1504.fifo_wr_block = 0;
    assign fifo_intf_1504.finish = finish;
    csv_file_dump fifo_csv_dumper_1504;
    csv_file_dump cstatus_csv_dumper_1504;
    df_fifo_monitor fifo_monitor_1504;
    df_fifo_intf fifo_intf_1505(clock,reset);
    assign fifo_intf_1505.rd_en = AESL_inst_myproject.layer3_out_152_U.if_read & AESL_inst_myproject.layer3_out_152_U.if_empty_n;
    assign fifo_intf_1505.wr_en = AESL_inst_myproject.layer3_out_152_U.if_write & AESL_inst_myproject.layer3_out_152_U.if_full_n;
    assign fifo_intf_1505.fifo_rd_block = 0;
    assign fifo_intf_1505.fifo_wr_block = 0;
    assign fifo_intf_1505.finish = finish;
    csv_file_dump fifo_csv_dumper_1505;
    csv_file_dump cstatus_csv_dumper_1505;
    df_fifo_monitor fifo_monitor_1505;
    df_fifo_intf fifo_intf_1506(clock,reset);
    assign fifo_intf_1506.rd_en = AESL_inst_myproject.layer3_out_153_U.if_read & AESL_inst_myproject.layer3_out_153_U.if_empty_n;
    assign fifo_intf_1506.wr_en = AESL_inst_myproject.layer3_out_153_U.if_write & AESL_inst_myproject.layer3_out_153_U.if_full_n;
    assign fifo_intf_1506.fifo_rd_block = 0;
    assign fifo_intf_1506.fifo_wr_block = 0;
    assign fifo_intf_1506.finish = finish;
    csv_file_dump fifo_csv_dumper_1506;
    csv_file_dump cstatus_csv_dumper_1506;
    df_fifo_monitor fifo_monitor_1506;
    df_fifo_intf fifo_intf_1507(clock,reset);
    assign fifo_intf_1507.rd_en = AESL_inst_myproject.layer3_out_154_U.if_read & AESL_inst_myproject.layer3_out_154_U.if_empty_n;
    assign fifo_intf_1507.wr_en = AESL_inst_myproject.layer3_out_154_U.if_write & AESL_inst_myproject.layer3_out_154_U.if_full_n;
    assign fifo_intf_1507.fifo_rd_block = 0;
    assign fifo_intf_1507.fifo_wr_block = 0;
    assign fifo_intf_1507.finish = finish;
    csv_file_dump fifo_csv_dumper_1507;
    csv_file_dump cstatus_csv_dumper_1507;
    df_fifo_monitor fifo_monitor_1507;
    df_fifo_intf fifo_intf_1508(clock,reset);
    assign fifo_intf_1508.rd_en = AESL_inst_myproject.layer3_out_155_U.if_read & AESL_inst_myproject.layer3_out_155_U.if_empty_n;
    assign fifo_intf_1508.wr_en = AESL_inst_myproject.layer3_out_155_U.if_write & AESL_inst_myproject.layer3_out_155_U.if_full_n;
    assign fifo_intf_1508.fifo_rd_block = 0;
    assign fifo_intf_1508.fifo_wr_block = 0;
    assign fifo_intf_1508.finish = finish;
    csv_file_dump fifo_csv_dumper_1508;
    csv_file_dump cstatus_csv_dumper_1508;
    df_fifo_monitor fifo_monitor_1508;
    df_fifo_intf fifo_intf_1509(clock,reset);
    assign fifo_intf_1509.rd_en = AESL_inst_myproject.layer3_out_156_U.if_read & AESL_inst_myproject.layer3_out_156_U.if_empty_n;
    assign fifo_intf_1509.wr_en = AESL_inst_myproject.layer3_out_156_U.if_write & AESL_inst_myproject.layer3_out_156_U.if_full_n;
    assign fifo_intf_1509.fifo_rd_block = 0;
    assign fifo_intf_1509.fifo_wr_block = 0;
    assign fifo_intf_1509.finish = finish;
    csv_file_dump fifo_csv_dumper_1509;
    csv_file_dump cstatus_csv_dumper_1509;
    df_fifo_monitor fifo_monitor_1509;
    df_fifo_intf fifo_intf_1510(clock,reset);
    assign fifo_intf_1510.rd_en = AESL_inst_myproject.layer3_out_157_U.if_read & AESL_inst_myproject.layer3_out_157_U.if_empty_n;
    assign fifo_intf_1510.wr_en = AESL_inst_myproject.layer3_out_157_U.if_write & AESL_inst_myproject.layer3_out_157_U.if_full_n;
    assign fifo_intf_1510.fifo_rd_block = 0;
    assign fifo_intf_1510.fifo_wr_block = 0;
    assign fifo_intf_1510.finish = finish;
    csv_file_dump fifo_csv_dumper_1510;
    csv_file_dump cstatus_csv_dumper_1510;
    df_fifo_monitor fifo_monitor_1510;
    df_fifo_intf fifo_intf_1511(clock,reset);
    assign fifo_intf_1511.rd_en = AESL_inst_myproject.layer3_out_158_U.if_read & AESL_inst_myproject.layer3_out_158_U.if_empty_n;
    assign fifo_intf_1511.wr_en = AESL_inst_myproject.layer3_out_158_U.if_write & AESL_inst_myproject.layer3_out_158_U.if_full_n;
    assign fifo_intf_1511.fifo_rd_block = 0;
    assign fifo_intf_1511.fifo_wr_block = 0;
    assign fifo_intf_1511.finish = finish;
    csv_file_dump fifo_csv_dumper_1511;
    csv_file_dump cstatus_csv_dumper_1511;
    df_fifo_monitor fifo_monitor_1511;
    df_fifo_intf fifo_intf_1512(clock,reset);
    assign fifo_intf_1512.rd_en = AESL_inst_myproject.layer3_out_159_U.if_read & AESL_inst_myproject.layer3_out_159_U.if_empty_n;
    assign fifo_intf_1512.wr_en = AESL_inst_myproject.layer3_out_159_U.if_write & AESL_inst_myproject.layer3_out_159_U.if_full_n;
    assign fifo_intf_1512.fifo_rd_block = 0;
    assign fifo_intf_1512.fifo_wr_block = 0;
    assign fifo_intf_1512.finish = finish;
    csv_file_dump fifo_csv_dumper_1512;
    csv_file_dump cstatus_csv_dumper_1512;
    df_fifo_monitor fifo_monitor_1512;
    df_fifo_intf fifo_intf_1513(clock,reset);
    assign fifo_intf_1513.rd_en = AESL_inst_myproject.layer3_out_160_U.if_read & AESL_inst_myproject.layer3_out_160_U.if_empty_n;
    assign fifo_intf_1513.wr_en = AESL_inst_myproject.layer3_out_160_U.if_write & AESL_inst_myproject.layer3_out_160_U.if_full_n;
    assign fifo_intf_1513.fifo_rd_block = 0;
    assign fifo_intf_1513.fifo_wr_block = 0;
    assign fifo_intf_1513.finish = finish;
    csv_file_dump fifo_csv_dumper_1513;
    csv_file_dump cstatus_csv_dumper_1513;
    df_fifo_monitor fifo_monitor_1513;
    df_fifo_intf fifo_intf_1514(clock,reset);
    assign fifo_intf_1514.rd_en = AESL_inst_myproject.layer3_out_161_U.if_read & AESL_inst_myproject.layer3_out_161_U.if_empty_n;
    assign fifo_intf_1514.wr_en = AESL_inst_myproject.layer3_out_161_U.if_write & AESL_inst_myproject.layer3_out_161_U.if_full_n;
    assign fifo_intf_1514.fifo_rd_block = 0;
    assign fifo_intf_1514.fifo_wr_block = 0;
    assign fifo_intf_1514.finish = finish;
    csv_file_dump fifo_csv_dumper_1514;
    csv_file_dump cstatus_csv_dumper_1514;
    df_fifo_monitor fifo_monitor_1514;
    df_fifo_intf fifo_intf_1515(clock,reset);
    assign fifo_intf_1515.rd_en = AESL_inst_myproject.layer3_out_162_U.if_read & AESL_inst_myproject.layer3_out_162_U.if_empty_n;
    assign fifo_intf_1515.wr_en = AESL_inst_myproject.layer3_out_162_U.if_write & AESL_inst_myproject.layer3_out_162_U.if_full_n;
    assign fifo_intf_1515.fifo_rd_block = 0;
    assign fifo_intf_1515.fifo_wr_block = 0;
    assign fifo_intf_1515.finish = finish;
    csv_file_dump fifo_csv_dumper_1515;
    csv_file_dump cstatus_csv_dumper_1515;
    df_fifo_monitor fifo_monitor_1515;
    df_fifo_intf fifo_intf_1516(clock,reset);
    assign fifo_intf_1516.rd_en = AESL_inst_myproject.layer3_out_163_U.if_read & AESL_inst_myproject.layer3_out_163_U.if_empty_n;
    assign fifo_intf_1516.wr_en = AESL_inst_myproject.layer3_out_163_U.if_write & AESL_inst_myproject.layer3_out_163_U.if_full_n;
    assign fifo_intf_1516.fifo_rd_block = 0;
    assign fifo_intf_1516.fifo_wr_block = 0;
    assign fifo_intf_1516.finish = finish;
    csv_file_dump fifo_csv_dumper_1516;
    csv_file_dump cstatus_csv_dumper_1516;
    df_fifo_monitor fifo_monitor_1516;
    df_fifo_intf fifo_intf_1517(clock,reset);
    assign fifo_intf_1517.rd_en = AESL_inst_myproject.layer3_out_164_U.if_read & AESL_inst_myproject.layer3_out_164_U.if_empty_n;
    assign fifo_intf_1517.wr_en = AESL_inst_myproject.layer3_out_164_U.if_write & AESL_inst_myproject.layer3_out_164_U.if_full_n;
    assign fifo_intf_1517.fifo_rd_block = 0;
    assign fifo_intf_1517.fifo_wr_block = 0;
    assign fifo_intf_1517.finish = finish;
    csv_file_dump fifo_csv_dumper_1517;
    csv_file_dump cstatus_csv_dumper_1517;
    df_fifo_monitor fifo_monitor_1517;
    df_fifo_intf fifo_intf_1518(clock,reset);
    assign fifo_intf_1518.rd_en = AESL_inst_myproject.layer3_out_165_U.if_read & AESL_inst_myproject.layer3_out_165_U.if_empty_n;
    assign fifo_intf_1518.wr_en = AESL_inst_myproject.layer3_out_165_U.if_write & AESL_inst_myproject.layer3_out_165_U.if_full_n;
    assign fifo_intf_1518.fifo_rd_block = 0;
    assign fifo_intf_1518.fifo_wr_block = 0;
    assign fifo_intf_1518.finish = finish;
    csv_file_dump fifo_csv_dumper_1518;
    csv_file_dump cstatus_csv_dumper_1518;
    df_fifo_monitor fifo_monitor_1518;
    df_fifo_intf fifo_intf_1519(clock,reset);
    assign fifo_intf_1519.rd_en = AESL_inst_myproject.layer3_out_166_U.if_read & AESL_inst_myproject.layer3_out_166_U.if_empty_n;
    assign fifo_intf_1519.wr_en = AESL_inst_myproject.layer3_out_166_U.if_write & AESL_inst_myproject.layer3_out_166_U.if_full_n;
    assign fifo_intf_1519.fifo_rd_block = 0;
    assign fifo_intf_1519.fifo_wr_block = 0;
    assign fifo_intf_1519.finish = finish;
    csv_file_dump fifo_csv_dumper_1519;
    csv_file_dump cstatus_csv_dumper_1519;
    df_fifo_monitor fifo_monitor_1519;
    df_fifo_intf fifo_intf_1520(clock,reset);
    assign fifo_intf_1520.rd_en = AESL_inst_myproject.layer3_out_167_U.if_read & AESL_inst_myproject.layer3_out_167_U.if_empty_n;
    assign fifo_intf_1520.wr_en = AESL_inst_myproject.layer3_out_167_U.if_write & AESL_inst_myproject.layer3_out_167_U.if_full_n;
    assign fifo_intf_1520.fifo_rd_block = 0;
    assign fifo_intf_1520.fifo_wr_block = 0;
    assign fifo_intf_1520.finish = finish;
    csv_file_dump fifo_csv_dumper_1520;
    csv_file_dump cstatus_csv_dumper_1520;
    df_fifo_monitor fifo_monitor_1520;
    df_fifo_intf fifo_intf_1521(clock,reset);
    assign fifo_intf_1521.rd_en = AESL_inst_myproject.layer3_out_168_U.if_read & AESL_inst_myproject.layer3_out_168_U.if_empty_n;
    assign fifo_intf_1521.wr_en = AESL_inst_myproject.layer3_out_168_U.if_write & AESL_inst_myproject.layer3_out_168_U.if_full_n;
    assign fifo_intf_1521.fifo_rd_block = 0;
    assign fifo_intf_1521.fifo_wr_block = 0;
    assign fifo_intf_1521.finish = finish;
    csv_file_dump fifo_csv_dumper_1521;
    csv_file_dump cstatus_csv_dumper_1521;
    df_fifo_monitor fifo_monitor_1521;
    df_fifo_intf fifo_intf_1522(clock,reset);
    assign fifo_intf_1522.rd_en = AESL_inst_myproject.layer3_out_169_U.if_read & AESL_inst_myproject.layer3_out_169_U.if_empty_n;
    assign fifo_intf_1522.wr_en = AESL_inst_myproject.layer3_out_169_U.if_write & AESL_inst_myproject.layer3_out_169_U.if_full_n;
    assign fifo_intf_1522.fifo_rd_block = 0;
    assign fifo_intf_1522.fifo_wr_block = 0;
    assign fifo_intf_1522.finish = finish;
    csv_file_dump fifo_csv_dumper_1522;
    csv_file_dump cstatus_csv_dumper_1522;
    df_fifo_monitor fifo_monitor_1522;
    df_fifo_intf fifo_intf_1523(clock,reset);
    assign fifo_intf_1523.rd_en = AESL_inst_myproject.layer3_out_170_U.if_read & AESL_inst_myproject.layer3_out_170_U.if_empty_n;
    assign fifo_intf_1523.wr_en = AESL_inst_myproject.layer3_out_170_U.if_write & AESL_inst_myproject.layer3_out_170_U.if_full_n;
    assign fifo_intf_1523.fifo_rd_block = 0;
    assign fifo_intf_1523.fifo_wr_block = 0;
    assign fifo_intf_1523.finish = finish;
    csv_file_dump fifo_csv_dumper_1523;
    csv_file_dump cstatus_csv_dumper_1523;
    df_fifo_monitor fifo_monitor_1523;
    df_fifo_intf fifo_intf_1524(clock,reset);
    assign fifo_intf_1524.rd_en = AESL_inst_myproject.layer3_out_171_U.if_read & AESL_inst_myproject.layer3_out_171_U.if_empty_n;
    assign fifo_intf_1524.wr_en = AESL_inst_myproject.layer3_out_171_U.if_write & AESL_inst_myproject.layer3_out_171_U.if_full_n;
    assign fifo_intf_1524.fifo_rd_block = 0;
    assign fifo_intf_1524.fifo_wr_block = 0;
    assign fifo_intf_1524.finish = finish;
    csv_file_dump fifo_csv_dumper_1524;
    csv_file_dump cstatus_csv_dumper_1524;
    df_fifo_monitor fifo_monitor_1524;
    df_fifo_intf fifo_intf_1525(clock,reset);
    assign fifo_intf_1525.rd_en = AESL_inst_myproject.layer3_out_172_U.if_read & AESL_inst_myproject.layer3_out_172_U.if_empty_n;
    assign fifo_intf_1525.wr_en = AESL_inst_myproject.layer3_out_172_U.if_write & AESL_inst_myproject.layer3_out_172_U.if_full_n;
    assign fifo_intf_1525.fifo_rd_block = 0;
    assign fifo_intf_1525.fifo_wr_block = 0;
    assign fifo_intf_1525.finish = finish;
    csv_file_dump fifo_csv_dumper_1525;
    csv_file_dump cstatus_csv_dumper_1525;
    df_fifo_monitor fifo_monitor_1525;
    df_fifo_intf fifo_intf_1526(clock,reset);
    assign fifo_intf_1526.rd_en = AESL_inst_myproject.layer3_out_173_U.if_read & AESL_inst_myproject.layer3_out_173_U.if_empty_n;
    assign fifo_intf_1526.wr_en = AESL_inst_myproject.layer3_out_173_U.if_write & AESL_inst_myproject.layer3_out_173_U.if_full_n;
    assign fifo_intf_1526.fifo_rd_block = 0;
    assign fifo_intf_1526.fifo_wr_block = 0;
    assign fifo_intf_1526.finish = finish;
    csv_file_dump fifo_csv_dumper_1526;
    csv_file_dump cstatus_csv_dumper_1526;
    df_fifo_monitor fifo_monitor_1526;
    df_fifo_intf fifo_intf_1527(clock,reset);
    assign fifo_intf_1527.rd_en = AESL_inst_myproject.layer3_out_174_U.if_read & AESL_inst_myproject.layer3_out_174_U.if_empty_n;
    assign fifo_intf_1527.wr_en = AESL_inst_myproject.layer3_out_174_U.if_write & AESL_inst_myproject.layer3_out_174_U.if_full_n;
    assign fifo_intf_1527.fifo_rd_block = 0;
    assign fifo_intf_1527.fifo_wr_block = 0;
    assign fifo_intf_1527.finish = finish;
    csv_file_dump fifo_csv_dumper_1527;
    csv_file_dump cstatus_csv_dumper_1527;
    df_fifo_monitor fifo_monitor_1527;
    df_fifo_intf fifo_intf_1528(clock,reset);
    assign fifo_intf_1528.rd_en = AESL_inst_myproject.layer3_out_175_U.if_read & AESL_inst_myproject.layer3_out_175_U.if_empty_n;
    assign fifo_intf_1528.wr_en = AESL_inst_myproject.layer3_out_175_U.if_write & AESL_inst_myproject.layer3_out_175_U.if_full_n;
    assign fifo_intf_1528.fifo_rd_block = 0;
    assign fifo_intf_1528.fifo_wr_block = 0;
    assign fifo_intf_1528.finish = finish;
    csv_file_dump fifo_csv_dumper_1528;
    csv_file_dump cstatus_csv_dumper_1528;
    df_fifo_monitor fifo_monitor_1528;
    df_fifo_intf fifo_intf_1529(clock,reset);
    assign fifo_intf_1529.rd_en = AESL_inst_myproject.layer3_out_176_U.if_read & AESL_inst_myproject.layer3_out_176_U.if_empty_n;
    assign fifo_intf_1529.wr_en = AESL_inst_myproject.layer3_out_176_U.if_write & AESL_inst_myproject.layer3_out_176_U.if_full_n;
    assign fifo_intf_1529.fifo_rd_block = 0;
    assign fifo_intf_1529.fifo_wr_block = 0;
    assign fifo_intf_1529.finish = finish;
    csv_file_dump fifo_csv_dumper_1529;
    csv_file_dump cstatus_csv_dumper_1529;
    df_fifo_monitor fifo_monitor_1529;
    df_fifo_intf fifo_intf_1530(clock,reset);
    assign fifo_intf_1530.rd_en = AESL_inst_myproject.layer3_out_177_U.if_read & AESL_inst_myproject.layer3_out_177_U.if_empty_n;
    assign fifo_intf_1530.wr_en = AESL_inst_myproject.layer3_out_177_U.if_write & AESL_inst_myproject.layer3_out_177_U.if_full_n;
    assign fifo_intf_1530.fifo_rd_block = 0;
    assign fifo_intf_1530.fifo_wr_block = 0;
    assign fifo_intf_1530.finish = finish;
    csv_file_dump fifo_csv_dumper_1530;
    csv_file_dump cstatus_csv_dumper_1530;
    df_fifo_monitor fifo_monitor_1530;
    df_fifo_intf fifo_intf_1531(clock,reset);
    assign fifo_intf_1531.rd_en = AESL_inst_myproject.layer3_out_178_U.if_read & AESL_inst_myproject.layer3_out_178_U.if_empty_n;
    assign fifo_intf_1531.wr_en = AESL_inst_myproject.layer3_out_178_U.if_write & AESL_inst_myproject.layer3_out_178_U.if_full_n;
    assign fifo_intf_1531.fifo_rd_block = 0;
    assign fifo_intf_1531.fifo_wr_block = 0;
    assign fifo_intf_1531.finish = finish;
    csv_file_dump fifo_csv_dumper_1531;
    csv_file_dump cstatus_csv_dumper_1531;
    df_fifo_monitor fifo_monitor_1531;
    df_fifo_intf fifo_intf_1532(clock,reset);
    assign fifo_intf_1532.rd_en = AESL_inst_myproject.layer3_out_179_U.if_read & AESL_inst_myproject.layer3_out_179_U.if_empty_n;
    assign fifo_intf_1532.wr_en = AESL_inst_myproject.layer3_out_179_U.if_write & AESL_inst_myproject.layer3_out_179_U.if_full_n;
    assign fifo_intf_1532.fifo_rd_block = 0;
    assign fifo_intf_1532.fifo_wr_block = 0;
    assign fifo_intf_1532.finish = finish;
    csv_file_dump fifo_csv_dumper_1532;
    csv_file_dump cstatus_csv_dumper_1532;
    df_fifo_monitor fifo_monitor_1532;
    df_fifo_intf fifo_intf_1533(clock,reset);
    assign fifo_intf_1533.rd_en = AESL_inst_myproject.layer3_out_180_U.if_read & AESL_inst_myproject.layer3_out_180_U.if_empty_n;
    assign fifo_intf_1533.wr_en = AESL_inst_myproject.layer3_out_180_U.if_write & AESL_inst_myproject.layer3_out_180_U.if_full_n;
    assign fifo_intf_1533.fifo_rd_block = 0;
    assign fifo_intf_1533.fifo_wr_block = 0;
    assign fifo_intf_1533.finish = finish;
    csv_file_dump fifo_csv_dumper_1533;
    csv_file_dump cstatus_csv_dumper_1533;
    df_fifo_monitor fifo_monitor_1533;
    df_fifo_intf fifo_intf_1534(clock,reset);
    assign fifo_intf_1534.rd_en = AESL_inst_myproject.layer3_out_181_U.if_read & AESL_inst_myproject.layer3_out_181_U.if_empty_n;
    assign fifo_intf_1534.wr_en = AESL_inst_myproject.layer3_out_181_U.if_write & AESL_inst_myproject.layer3_out_181_U.if_full_n;
    assign fifo_intf_1534.fifo_rd_block = 0;
    assign fifo_intf_1534.fifo_wr_block = 0;
    assign fifo_intf_1534.finish = finish;
    csv_file_dump fifo_csv_dumper_1534;
    csv_file_dump cstatus_csv_dumper_1534;
    df_fifo_monitor fifo_monitor_1534;
    df_fifo_intf fifo_intf_1535(clock,reset);
    assign fifo_intf_1535.rd_en = AESL_inst_myproject.layer3_out_182_U.if_read & AESL_inst_myproject.layer3_out_182_U.if_empty_n;
    assign fifo_intf_1535.wr_en = AESL_inst_myproject.layer3_out_182_U.if_write & AESL_inst_myproject.layer3_out_182_U.if_full_n;
    assign fifo_intf_1535.fifo_rd_block = 0;
    assign fifo_intf_1535.fifo_wr_block = 0;
    assign fifo_intf_1535.finish = finish;
    csv_file_dump fifo_csv_dumper_1535;
    csv_file_dump cstatus_csv_dumper_1535;
    df_fifo_monitor fifo_monitor_1535;
    df_fifo_intf fifo_intf_1536(clock,reset);
    assign fifo_intf_1536.rd_en = AESL_inst_myproject.layer3_out_183_U.if_read & AESL_inst_myproject.layer3_out_183_U.if_empty_n;
    assign fifo_intf_1536.wr_en = AESL_inst_myproject.layer3_out_183_U.if_write & AESL_inst_myproject.layer3_out_183_U.if_full_n;
    assign fifo_intf_1536.fifo_rd_block = 0;
    assign fifo_intf_1536.fifo_wr_block = 0;
    assign fifo_intf_1536.finish = finish;
    csv_file_dump fifo_csv_dumper_1536;
    csv_file_dump cstatus_csv_dumper_1536;
    df_fifo_monitor fifo_monitor_1536;
    df_fifo_intf fifo_intf_1537(clock,reset);
    assign fifo_intf_1537.rd_en = AESL_inst_myproject.layer3_out_184_U.if_read & AESL_inst_myproject.layer3_out_184_U.if_empty_n;
    assign fifo_intf_1537.wr_en = AESL_inst_myproject.layer3_out_184_U.if_write & AESL_inst_myproject.layer3_out_184_U.if_full_n;
    assign fifo_intf_1537.fifo_rd_block = 0;
    assign fifo_intf_1537.fifo_wr_block = 0;
    assign fifo_intf_1537.finish = finish;
    csv_file_dump fifo_csv_dumper_1537;
    csv_file_dump cstatus_csv_dumper_1537;
    df_fifo_monitor fifo_monitor_1537;
    df_fifo_intf fifo_intf_1538(clock,reset);
    assign fifo_intf_1538.rd_en = AESL_inst_myproject.layer3_out_185_U.if_read & AESL_inst_myproject.layer3_out_185_U.if_empty_n;
    assign fifo_intf_1538.wr_en = AESL_inst_myproject.layer3_out_185_U.if_write & AESL_inst_myproject.layer3_out_185_U.if_full_n;
    assign fifo_intf_1538.fifo_rd_block = 0;
    assign fifo_intf_1538.fifo_wr_block = 0;
    assign fifo_intf_1538.finish = finish;
    csv_file_dump fifo_csv_dumper_1538;
    csv_file_dump cstatus_csv_dumper_1538;
    df_fifo_monitor fifo_monitor_1538;
    df_fifo_intf fifo_intf_1539(clock,reset);
    assign fifo_intf_1539.rd_en = AESL_inst_myproject.layer3_out_186_U.if_read & AESL_inst_myproject.layer3_out_186_U.if_empty_n;
    assign fifo_intf_1539.wr_en = AESL_inst_myproject.layer3_out_186_U.if_write & AESL_inst_myproject.layer3_out_186_U.if_full_n;
    assign fifo_intf_1539.fifo_rd_block = 0;
    assign fifo_intf_1539.fifo_wr_block = 0;
    assign fifo_intf_1539.finish = finish;
    csv_file_dump fifo_csv_dumper_1539;
    csv_file_dump cstatus_csv_dumper_1539;
    df_fifo_monitor fifo_monitor_1539;
    df_fifo_intf fifo_intf_1540(clock,reset);
    assign fifo_intf_1540.rd_en = AESL_inst_myproject.layer3_out_187_U.if_read & AESL_inst_myproject.layer3_out_187_U.if_empty_n;
    assign fifo_intf_1540.wr_en = AESL_inst_myproject.layer3_out_187_U.if_write & AESL_inst_myproject.layer3_out_187_U.if_full_n;
    assign fifo_intf_1540.fifo_rd_block = 0;
    assign fifo_intf_1540.fifo_wr_block = 0;
    assign fifo_intf_1540.finish = finish;
    csv_file_dump fifo_csv_dumper_1540;
    csv_file_dump cstatus_csv_dumper_1540;
    df_fifo_monitor fifo_monitor_1540;
    df_fifo_intf fifo_intf_1541(clock,reset);
    assign fifo_intf_1541.rd_en = AESL_inst_myproject.layer3_out_188_U.if_read & AESL_inst_myproject.layer3_out_188_U.if_empty_n;
    assign fifo_intf_1541.wr_en = AESL_inst_myproject.layer3_out_188_U.if_write & AESL_inst_myproject.layer3_out_188_U.if_full_n;
    assign fifo_intf_1541.fifo_rd_block = 0;
    assign fifo_intf_1541.fifo_wr_block = 0;
    assign fifo_intf_1541.finish = finish;
    csv_file_dump fifo_csv_dumper_1541;
    csv_file_dump cstatus_csv_dumper_1541;
    df_fifo_monitor fifo_monitor_1541;
    df_fifo_intf fifo_intf_1542(clock,reset);
    assign fifo_intf_1542.rd_en = AESL_inst_myproject.layer3_out_189_U.if_read & AESL_inst_myproject.layer3_out_189_U.if_empty_n;
    assign fifo_intf_1542.wr_en = AESL_inst_myproject.layer3_out_189_U.if_write & AESL_inst_myproject.layer3_out_189_U.if_full_n;
    assign fifo_intf_1542.fifo_rd_block = 0;
    assign fifo_intf_1542.fifo_wr_block = 0;
    assign fifo_intf_1542.finish = finish;
    csv_file_dump fifo_csv_dumper_1542;
    csv_file_dump cstatus_csv_dumper_1542;
    df_fifo_monitor fifo_monitor_1542;
    df_fifo_intf fifo_intf_1543(clock,reset);
    assign fifo_intf_1543.rd_en = AESL_inst_myproject.layer3_out_190_U.if_read & AESL_inst_myproject.layer3_out_190_U.if_empty_n;
    assign fifo_intf_1543.wr_en = AESL_inst_myproject.layer3_out_190_U.if_write & AESL_inst_myproject.layer3_out_190_U.if_full_n;
    assign fifo_intf_1543.fifo_rd_block = 0;
    assign fifo_intf_1543.fifo_wr_block = 0;
    assign fifo_intf_1543.finish = finish;
    csv_file_dump fifo_csv_dumper_1543;
    csv_file_dump cstatus_csv_dumper_1543;
    df_fifo_monitor fifo_monitor_1543;
    df_fifo_intf fifo_intf_1544(clock,reset);
    assign fifo_intf_1544.rd_en = AESL_inst_myproject.layer3_out_191_U.if_read & AESL_inst_myproject.layer3_out_191_U.if_empty_n;
    assign fifo_intf_1544.wr_en = AESL_inst_myproject.layer3_out_191_U.if_write & AESL_inst_myproject.layer3_out_191_U.if_full_n;
    assign fifo_intf_1544.fifo_rd_block = 0;
    assign fifo_intf_1544.fifo_wr_block = 0;
    assign fifo_intf_1544.finish = finish;
    csv_file_dump fifo_csv_dumper_1544;
    csv_file_dump cstatus_csv_dumper_1544;
    df_fifo_monitor fifo_monitor_1544;
    df_fifo_intf fifo_intf_1545(clock,reset);
    assign fifo_intf_1545.rd_en = AESL_inst_myproject.layer3_out_192_U.if_read & AESL_inst_myproject.layer3_out_192_U.if_empty_n;
    assign fifo_intf_1545.wr_en = AESL_inst_myproject.layer3_out_192_U.if_write & AESL_inst_myproject.layer3_out_192_U.if_full_n;
    assign fifo_intf_1545.fifo_rd_block = 0;
    assign fifo_intf_1545.fifo_wr_block = 0;
    assign fifo_intf_1545.finish = finish;
    csv_file_dump fifo_csv_dumper_1545;
    csv_file_dump cstatus_csv_dumper_1545;
    df_fifo_monitor fifo_monitor_1545;
    df_fifo_intf fifo_intf_1546(clock,reset);
    assign fifo_intf_1546.rd_en = AESL_inst_myproject.layer3_out_193_U.if_read & AESL_inst_myproject.layer3_out_193_U.if_empty_n;
    assign fifo_intf_1546.wr_en = AESL_inst_myproject.layer3_out_193_U.if_write & AESL_inst_myproject.layer3_out_193_U.if_full_n;
    assign fifo_intf_1546.fifo_rd_block = 0;
    assign fifo_intf_1546.fifo_wr_block = 0;
    assign fifo_intf_1546.finish = finish;
    csv_file_dump fifo_csv_dumper_1546;
    csv_file_dump cstatus_csv_dumper_1546;
    df_fifo_monitor fifo_monitor_1546;
    df_fifo_intf fifo_intf_1547(clock,reset);
    assign fifo_intf_1547.rd_en = AESL_inst_myproject.layer3_out_194_U.if_read & AESL_inst_myproject.layer3_out_194_U.if_empty_n;
    assign fifo_intf_1547.wr_en = AESL_inst_myproject.layer3_out_194_U.if_write & AESL_inst_myproject.layer3_out_194_U.if_full_n;
    assign fifo_intf_1547.fifo_rd_block = 0;
    assign fifo_intf_1547.fifo_wr_block = 0;
    assign fifo_intf_1547.finish = finish;
    csv_file_dump fifo_csv_dumper_1547;
    csv_file_dump cstatus_csv_dumper_1547;
    df_fifo_monitor fifo_monitor_1547;
    df_fifo_intf fifo_intf_1548(clock,reset);
    assign fifo_intf_1548.rd_en = AESL_inst_myproject.layer3_out_195_U.if_read & AESL_inst_myproject.layer3_out_195_U.if_empty_n;
    assign fifo_intf_1548.wr_en = AESL_inst_myproject.layer3_out_195_U.if_write & AESL_inst_myproject.layer3_out_195_U.if_full_n;
    assign fifo_intf_1548.fifo_rd_block = 0;
    assign fifo_intf_1548.fifo_wr_block = 0;
    assign fifo_intf_1548.finish = finish;
    csv_file_dump fifo_csv_dumper_1548;
    csv_file_dump cstatus_csv_dumper_1548;
    df_fifo_monitor fifo_monitor_1548;
    df_fifo_intf fifo_intf_1549(clock,reset);
    assign fifo_intf_1549.rd_en = AESL_inst_myproject.layer3_out_196_U.if_read & AESL_inst_myproject.layer3_out_196_U.if_empty_n;
    assign fifo_intf_1549.wr_en = AESL_inst_myproject.layer3_out_196_U.if_write & AESL_inst_myproject.layer3_out_196_U.if_full_n;
    assign fifo_intf_1549.fifo_rd_block = 0;
    assign fifo_intf_1549.fifo_wr_block = 0;
    assign fifo_intf_1549.finish = finish;
    csv_file_dump fifo_csv_dumper_1549;
    csv_file_dump cstatus_csv_dumper_1549;
    df_fifo_monitor fifo_monitor_1549;
    df_fifo_intf fifo_intf_1550(clock,reset);
    assign fifo_intf_1550.rd_en = AESL_inst_myproject.layer3_out_197_U.if_read & AESL_inst_myproject.layer3_out_197_U.if_empty_n;
    assign fifo_intf_1550.wr_en = AESL_inst_myproject.layer3_out_197_U.if_write & AESL_inst_myproject.layer3_out_197_U.if_full_n;
    assign fifo_intf_1550.fifo_rd_block = 0;
    assign fifo_intf_1550.fifo_wr_block = 0;
    assign fifo_intf_1550.finish = finish;
    csv_file_dump fifo_csv_dumper_1550;
    csv_file_dump cstatus_csv_dumper_1550;
    df_fifo_monitor fifo_monitor_1550;
    df_fifo_intf fifo_intf_1551(clock,reset);
    assign fifo_intf_1551.rd_en = AESL_inst_myproject.layer3_out_198_U.if_read & AESL_inst_myproject.layer3_out_198_U.if_empty_n;
    assign fifo_intf_1551.wr_en = AESL_inst_myproject.layer3_out_198_U.if_write & AESL_inst_myproject.layer3_out_198_U.if_full_n;
    assign fifo_intf_1551.fifo_rd_block = 0;
    assign fifo_intf_1551.fifo_wr_block = 0;
    assign fifo_intf_1551.finish = finish;
    csv_file_dump fifo_csv_dumper_1551;
    csv_file_dump cstatus_csv_dumper_1551;
    df_fifo_monitor fifo_monitor_1551;
    df_fifo_intf fifo_intf_1552(clock,reset);
    assign fifo_intf_1552.rd_en = AESL_inst_myproject.layer3_out_199_U.if_read & AESL_inst_myproject.layer3_out_199_U.if_empty_n;
    assign fifo_intf_1552.wr_en = AESL_inst_myproject.layer3_out_199_U.if_write & AESL_inst_myproject.layer3_out_199_U.if_full_n;
    assign fifo_intf_1552.fifo_rd_block = 0;
    assign fifo_intf_1552.fifo_wr_block = 0;
    assign fifo_intf_1552.finish = finish;
    csv_file_dump fifo_csv_dumper_1552;
    csv_file_dump cstatus_csv_dumper_1552;
    df_fifo_monitor fifo_monitor_1552;
    df_fifo_intf fifo_intf_1553(clock,reset);
    assign fifo_intf_1553.rd_en = AESL_inst_myproject.layer3_out_200_U.if_read & AESL_inst_myproject.layer3_out_200_U.if_empty_n;
    assign fifo_intf_1553.wr_en = AESL_inst_myproject.layer3_out_200_U.if_write & AESL_inst_myproject.layer3_out_200_U.if_full_n;
    assign fifo_intf_1553.fifo_rd_block = 0;
    assign fifo_intf_1553.fifo_wr_block = 0;
    assign fifo_intf_1553.finish = finish;
    csv_file_dump fifo_csv_dumper_1553;
    csv_file_dump cstatus_csv_dumper_1553;
    df_fifo_monitor fifo_monitor_1553;
    df_fifo_intf fifo_intf_1554(clock,reset);
    assign fifo_intf_1554.rd_en = AESL_inst_myproject.layer3_out_201_U.if_read & AESL_inst_myproject.layer3_out_201_U.if_empty_n;
    assign fifo_intf_1554.wr_en = AESL_inst_myproject.layer3_out_201_U.if_write & AESL_inst_myproject.layer3_out_201_U.if_full_n;
    assign fifo_intf_1554.fifo_rd_block = 0;
    assign fifo_intf_1554.fifo_wr_block = 0;
    assign fifo_intf_1554.finish = finish;
    csv_file_dump fifo_csv_dumper_1554;
    csv_file_dump cstatus_csv_dumper_1554;
    df_fifo_monitor fifo_monitor_1554;
    df_fifo_intf fifo_intf_1555(clock,reset);
    assign fifo_intf_1555.rd_en = AESL_inst_myproject.layer3_out_202_U.if_read & AESL_inst_myproject.layer3_out_202_U.if_empty_n;
    assign fifo_intf_1555.wr_en = AESL_inst_myproject.layer3_out_202_U.if_write & AESL_inst_myproject.layer3_out_202_U.if_full_n;
    assign fifo_intf_1555.fifo_rd_block = 0;
    assign fifo_intf_1555.fifo_wr_block = 0;
    assign fifo_intf_1555.finish = finish;
    csv_file_dump fifo_csv_dumper_1555;
    csv_file_dump cstatus_csv_dumper_1555;
    df_fifo_monitor fifo_monitor_1555;
    df_fifo_intf fifo_intf_1556(clock,reset);
    assign fifo_intf_1556.rd_en = AESL_inst_myproject.layer3_out_203_U.if_read & AESL_inst_myproject.layer3_out_203_U.if_empty_n;
    assign fifo_intf_1556.wr_en = AESL_inst_myproject.layer3_out_203_U.if_write & AESL_inst_myproject.layer3_out_203_U.if_full_n;
    assign fifo_intf_1556.fifo_rd_block = 0;
    assign fifo_intf_1556.fifo_wr_block = 0;
    assign fifo_intf_1556.finish = finish;
    csv_file_dump fifo_csv_dumper_1556;
    csv_file_dump cstatus_csv_dumper_1556;
    df_fifo_monitor fifo_monitor_1556;
    df_fifo_intf fifo_intf_1557(clock,reset);
    assign fifo_intf_1557.rd_en = AESL_inst_myproject.layer3_out_204_U.if_read & AESL_inst_myproject.layer3_out_204_U.if_empty_n;
    assign fifo_intf_1557.wr_en = AESL_inst_myproject.layer3_out_204_U.if_write & AESL_inst_myproject.layer3_out_204_U.if_full_n;
    assign fifo_intf_1557.fifo_rd_block = 0;
    assign fifo_intf_1557.fifo_wr_block = 0;
    assign fifo_intf_1557.finish = finish;
    csv_file_dump fifo_csv_dumper_1557;
    csv_file_dump cstatus_csv_dumper_1557;
    df_fifo_monitor fifo_monitor_1557;
    df_fifo_intf fifo_intf_1558(clock,reset);
    assign fifo_intf_1558.rd_en = AESL_inst_myproject.layer3_out_205_U.if_read & AESL_inst_myproject.layer3_out_205_U.if_empty_n;
    assign fifo_intf_1558.wr_en = AESL_inst_myproject.layer3_out_205_U.if_write & AESL_inst_myproject.layer3_out_205_U.if_full_n;
    assign fifo_intf_1558.fifo_rd_block = 0;
    assign fifo_intf_1558.fifo_wr_block = 0;
    assign fifo_intf_1558.finish = finish;
    csv_file_dump fifo_csv_dumper_1558;
    csv_file_dump cstatus_csv_dumper_1558;
    df_fifo_monitor fifo_monitor_1558;
    df_fifo_intf fifo_intf_1559(clock,reset);
    assign fifo_intf_1559.rd_en = AESL_inst_myproject.layer3_out_206_U.if_read & AESL_inst_myproject.layer3_out_206_U.if_empty_n;
    assign fifo_intf_1559.wr_en = AESL_inst_myproject.layer3_out_206_U.if_write & AESL_inst_myproject.layer3_out_206_U.if_full_n;
    assign fifo_intf_1559.fifo_rd_block = 0;
    assign fifo_intf_1559.fifo_wr_block = 0;
    assign fifo_intf_1559.finish = finish;
    csv_file_dump fifo_csv_dumper_1559;
    csv_file_dump cstatus_csv_dumper_1559;
    df_fifo_monitor fifo_monitor_1559;
    df_fifo_intf fifo_intf_1560(clock,reset);
    assign fifo_intf_1560.rd_en = AESL_inst_myproject.layer3_out_207_U.if_read & AESL_inst_myproject.layer3_out_207_U.if_empty_n;
    assign fifo_intf_1560.wr_en = AESL_inst_myproject.layer3_out_207_U.if_write & AESL_inst_myproject.layer3_out_207_U.if_full_n;
    assign fifo_intf_1560.fifo_rd_block = 0;
    assign fifo_intf_1560.fifo_wr_block = 0;
    assign fifo_intf_1560.finish = finish;
    csv_file_dump fifo_csv_dumper_1560;
    csv_file_dump cstatus_csv_dumper_1560;
    df_fifo_monitor fifo_monitor_1560;
    df_fifo_intf fifo_intf_1561(clock,reset);
    assign fifo_intf_1561.rd_en = AESL_inst_myproject.layer3_out_208_U.if_read & AESL_inst_myproject.layer3_out_208_U.if_empty_n;
    assign fifo_intf_1561.wr_en = AESL_inst_myproject.layer3_out_208_U.if_write & AESL_inst_myproject.layer3_out_208_U.if_full_n;
    assign fifo_intf_1561.fifo_rd_block = 0;
    assign fifo_intf_1561.fifo_wr_block = 0;
    assign fifo_intf_1561.finish = finish;
    csv_file_dump fifo_csv_dumper_1561;
    csv_file_dump cstatus_csv_dumper_1561;
    df_fifo_monitor fifo_monitor_1561;
    df_fifo_intf fifo_intf_1562(clock,reset);
    assign fifo_intf_1562.rd_en = AESL_inst_myproject.layer3_out_209_U.if_read & AESL_inst_myproject.layer3_out_209_U.if_empty_n;
    assign fifo_intf_1562.wr_en = AESL_inst_myproject.layer3_out_209_U.if_write & AESL_inst_myproject.layer3_out_209_U.if_full_n;
    assign fifo_intf_1562.fifo_rd_block = 0;
    assign fifo_intf_1562.fifo_wr_block = 0;
    assign fifo_intf_1562.finish = finish;
    csv_file_dump fifo_csv_dumper_1562;
    csv_file_dump cstatus_csv_dumper_1562;
    df_fifo_monitor fifo_monitor_1562;
    df_fifo_intf fifo_intf_1563(clock,reset);
    assign fifo_intf_1563.rd_en = AESL_inst_myproject.layer3_out_210_U.if_read & AESL_inst_myproject.layer3_out_210_U.if_empty_n;
    assign fifo_intf_1563.wr_en = AESL_inst_myproject.layer3_out_210_U.if_write & AESL_inst_myproject.layer3_out_210_U.if_full_n;
    assign fifo_intf_1563.fifo_rd_block = 0;
    assign fifo_intf_1563.fifo_wr_block = 0;
    assign fifo_intf_1563.finish = finish;
    csv_file_dump fifo_csv_dumper_1563;
    csv_file_dump cstatus_csv_dumper_1563;
    df_fifo_monitor fifo_monitor_1563;
    df_fifo_intf fifo_intf_1564(clock,reset);
    assign fifo_intf_1564.rd_en = AESL_inst_myproject.layer3_out_211_U.if_read & AESL_inst_myproject.layer3_out_211_U.if_empty_n;
    assign fifo_intf_1564.wr_en = AESL_inst_myproject.layer3_out_211_U.if_write & AESL_inst_myproject.layer3_out_211_U.if_full_n;
    assign fifo_intf_1564.fifo_rd_block = 0;
    assign fifo_intf_1564.fifo_wr_block = 0;
    assign fifo_intf_1564.finish = finish;
    csv_file_dump fifo_csv_dumper_1564;
    csv_file_dump cstatus_csv_dumper_1564;
    df_fifo_monitor fifo_monitor_1564;
    df_fifo_intf fifo_intf_1565(clock,reset);
    assign fifo_intf_1565.rd_en = AESL_inst_myproject.layer3_out_212_U.if_read & AESL_inst_myproject.layer3_out_212_U.if_empty_n;
    assign fifo_intf_1565.wr_en = AESL_inst_myproject.layer3_out_212_U.if_write & AESL_inst_myproject.layer3_out_212_U.if_full_n;
    assign fifo_intf_1565.fifo_rd_block = 0;
    assign fifo_intf_1565.fifo_wr_block = 0;
    assign fifo_intf_1565.finish = finish;
    csv_file_dump fifo_csv_dumper_1565;
    csv_file_dump cstatus_csv_dumper_1565;
    df_fifo_monitor fifo_monitor_1565;
    df_fifo_intf fifo_intf_1566(clock,reset);
    assign fifo_intf_1566.rd_en = AESL_inst_myproject.layer3_out_213_U.if_read & AESL_inst_myproject.layer3_out_213_U.if_empty_n;
    assign fifo_intf_1566.wr_en = AESL_inst_myproject.layer3_out_213_U.if_write & AESL_inst_myproject.layer3_out_213_U.if_full_n;
    assign fifo_intf_1566.fifo_rd_block = 0;
    assign fifo_intf_1566.fifo_wr_block = 0;
    assign fifo_intf_1566.finish = finish;
    csv_file_dump fifo_csv_dumper_1566;
    csv_file_dump cstatus_csv_dumper_1566;
    df_fifo_monitor fifo_monitor_1566;
    df_fifo_intf fifo_intf_1567(clock,reset);
    assign fifo_intf_1567.rd_en = AESL_inst_myproject.layer3_out_214_U.if_read & AESL_inst_myproject.layer3_out_214_U.if_empty_n;
    assign fifo_intf_1567.wr_en = AESL_inst_myproject.layer3_out_214_U.if_write & AESL_inst_myproject.layer3_out_214_U.if_full_n;
    assign fifo_intf_1567.fifo_rd_block = 0;
    assign fifo_intf_1567.fifo_wr_block = 0;
    assign fifo_intf_1567.finish = finish;
    csv_file_dump fifo_csv_dumper_1567;
    csv_file_dump cstatus_csv_dumper_1567;
    df_fifo_monitor fifo_monitor_1567;
    df_fifo_intf fifo_intf_1568(clock,reset);
    assign fifo_intf_1568.rd_en = AESL_inst_myproject.layer3_out_215_U.if_read & AESL_inst_myproject.layer3_out_215_U.if_empty_n;
    assign fifo_intf_1568.wr_en = AESL_inst_myproject.layer3_out_215_U.if_write & AESL_inst_myproject.layer3_out_215_U.if_full_n;
    assign fifo_intf_1568.fifo_rd_block = 0;
    assign fifo_intf_1568.fifo_wr_block = 0;
    assign fifo_intf_1568.finish = finish;
    csv_file_dump fifo_csv_dumper_1568;
    csv_file_dump cstatus_csv_dumper_1568;
    df_fifo_monitor fifo_monitor_1568;
    df_fifo_intf fifo_intf_1569(clock,reset);
    assign fifo_intf_1569.rd_en = AESL_inst_myproject.layer3_out_216_U.if_read & AESL_inst_myproject.layer3_out_216_U.if_empty_n;
    assign fifo_intf_1569.wr_en = AESL_inst_myproject.layer3_out_216_U.if_write & AESL_inst_myproject.layer3_out_216_U.if_full_n;
    assign fifo_intf_1569.fifo_rd_block = 0;
    assign fifo_intf_1569.fifo_wr_block = 0;
    assign fifo_intf_1569.finish = finish;
    csv_file_dump fifo_csv_dumper_1569;
    csv_file_dump cstatus_csv_dumper_1569;
    df_fifo_monitor fifo_monitor_1569;
    df_fifo_intf fifo_intf_1570(clock,reset);
    assign fifo_intf_1570.rd_en = AESL_inst_myproject.layer3_out_217_U.if_read & AESL_inst_myproject.layer3_out_217_U.if_empty_n;
    assign fifo_intf_1570.wr_en = AESL_inst_myproject.layer3_out_217_U.if_write & AESL_inst_myproject.layer3_out_217_U.if_full_n;
    assign fifo_intf_1570.fifo_rd_block = 0;
    assign fifo_intf_1570.fifo_wr_block = 0;
    assign fifo_intf_1570.finish = finish;
    csv_file_dump fifo_csv_dumper_1570;
    csv_file_dump cstatus_csv_dumper_1570;
    df_fifo_monitor fifo_monitor_1570;
    df_fifo_intf fifo_intf_1571(clock,reset);
    assign fifo_intf_1571.rd_en = AESL_inst_myproject.layer3_out_218_U.if_read & AESL_inst_myproject.layer3_out_218_U.if_empty_n;
    assign fifo_intf_1571.wr_en = AESL_inst_myproject.layer3_out_218_U.if_write & AESL_inst_myproject.layer3_out_218_U.if_full_n;
    assign fifo_intf_1571.fifo_rd_block = 0;
    assign fifo_intf_1571.fifo_wr_block = 0;
    assign fifo_intf_1571.finish = finish;
    csv_file_dump fifo_csv_dumper_1571;
    csv_file_dump cstatus_csv_dumper_1571;
    df_fifo_monitor fifo_monitor_1571;
    df_fifo_intf fifo_intf_1572(clock,reset);
    assign fifo_intf_1572.rd_en = AESL_inst_myproject.layer3_out_219_U.if_read & AESL_inst_myproject.layer3_out_219_U.if_empty_n;
    assign fifo_intf_1572.wr_en = AESL_inst_myproject.layer3_out_219_U.if_write & AESL_inst_myproject.layer3_out_219_U.if_full_n;
    assign fifo_intf_1572.fifo_rd_block = 0;
    assign fifo_intf_1572.fifo_wr_block = 0;
    assign fifo_intf_1572.finish = finish;
    csv_file_dump fifo_csv_dumper_1572;
    csv_file_dump cstatus_csv_dumper_1572;
    df_fifo_monitor fifo_monitor_1572;
    df_fifo_intf fifo_intf_1573(clock,reset);
    assign fifo_intf_1573.rd_en = AESL_inst_myproject.layer3_out_220_U.if_read & AESL_inst_myproject.layer3_out_220_U.if_empty_n;
    assign fifo_intf_1573.wr_en = AESL_inst_myproject.layer3_out_220_U.if_write & AESL_inst_myproject.layer3_out_220_U.if_full_n;
    assign fifo_intf_1573.fifo_rd_block = 0;
    assign fifo_intf_1573.fifo_wr_block = 0;
    assign fifo_intf_1573.finish = finish;
    csv_file_dump fifo_csv_dumper_1573;
    csv_file_dump cstatus_csv_dumper_1573;
    df_fifo_monitor fifo_monitor_1573;
    df_fifo_intf fifo_intf_1574(clock,reset);
    assign fifo_intf_1574.rd_en = AESL_inst_myproject.layer3_out_221_U.if_read & AESL_inst_myproject.layer3_out_221_U.if_empty_n;
    assign fifo_intf_1574.wr_en = AESL_inst_myproject.layer3_out_221_U.if_write & AESL_inst_myproject.layer3_out_221_U.if_full_n;
    assign fifo_intf_1574.fifo_rd_block = 0;
    assign fifo_intf_1574.fifo_wr_block = 0;
    assign fifo_intf_1574.finish = finish;
    csv_file_dump fifo_csv_dumper_1574;
    csv_file_dump cstatus_csv_dumper_1574;
    df_fifo_monitor fifo_monitor_1574;
    df_fifo_intf fifo_intf_1575(clock,reset);
    assign fifo_intf_1575.rd_en = AESL_inst_myproject.layer3_out_222_U.if_read & AESL_inst_myproject.layer3_out_222_U.if_empty_n;
    assign fifo_intf_1575.wr_en = AESL_inst_myproject.layer3_out_222_U.if_write & AESL_inst_myproject.layer3_out_222_U.if_full_n;
    assign fifo_intf_1575.fifo_rd_block = 0;
    assign fifo_intf_1575.fifo_wr_block = 0;
    assign fifo_intf_1575.finish = finish;
    csv_file_dump fifo_csv_dumper_1575;
    csv_file_dump cstatus_csv_dumper_1575;
    df_fifo_monitor fifo_monitor_1575;
    df_fifo_intf fifo_intf_1576(clock,reset);
    assign fifo_intf_1576.rd_en = AESL_inst_myproject.layer3_out_223_U.if_read & AESL_inst_myproject.layer3_out_223_U.if_empty_n;
    assign fifo_intf_1576.wr_en = AESL_inst_myproject.layer3_out_223_U.if_write & AESL_inst_myproject.layer3_out_223_U.if_full_n;
    assign fifo_intf_1576.fifo_rd_block = 0;
    assign fifo_intf_1576.fifo_wr_block = 0;
    assign fifo_intf_1576.finish = finish;
    csv_file_dump fifo_csv_dumper_1576;
    csv_file_dump cstatus_csv_dumper_1576;
    df_fifo_monitor fifo_monitor_1576;
    df_fifo_intf fifo_intf_1577(clock,reset);
    assign fifo_intf_1577.rd_en = AESL_inst_myproject.layer3_out_224_U.if_read & AESL_inst_myproject.layer3_out_224_U.if_empty_n;
    assign fifo_intf_1577.wr_en = AESL_inst_myproject.layer3_out_224_U.if_write & AESL_inst_myproject.layer3_out_224_U.if_full_n;
    assign fifo_intf_1577.fifo_rd_block = 0;
    assign fifo_intf_1577.fifo_wr_block = 0;
    assign fifo_intf_1577.finish = finish;
    csv_file_dump fifo_csv_dumper_1577;
    csv_file_dump cstatus_csv_dumper_1577;
    df_fifo_monitor fifo_monitor_1577;
    df_fifo_intf fifo_intf_1578(clock,reset);
    assign fifo_intf_1578.rd_en = AESL_inst_myproject.layer3_out_225_U.if_read & AESL_inst_myproject.layer3_out_225_U.if_empty_n;
    assign fifo_intf_1578.wr_en = AESL_inst_myproject.layer3_out_225_U.if_write & AESL_inst_myproject.layer3_out_225_U.if_full_n;
    assign fifo_intf_1578.fifo_rd_block = 0;
    assign fifo_intf_1578.fifo_wr_block = 0;
    assign fifo_intf_1578.finish = finish;
    csv_file_dump fifo_csv_dumper_1578;
    csv_file_dump cstatus_csv_dumper_1578;
    df_fifo_monitor fifo_monitor_1578;
    df_fifo_intf fifo_intf_1579(clock,reset);
    assign fifo_intf_1579.rd_en = AESL_inst_myproject.layer3_out_226_U.if_read & AESL_inst_myproject.layer3_out_226_U.if_empty_n;
    assign fifo_intf_1579.wr_en = AESL_inst_myproject.layer3_out_226_U.if_write & AESL_inst_myproject.layer3_out_226_U.if_full_n;
    assign fifo_intf_1579.fifo_rd_block = 0;
    assign fifo_intf_1579.fifo_wr_block = 0;
    assign fifo_intf_1579.finish = finish;
    csv_file_dump fifo_csv_dumper_1579;
    csv_file_dump cstatus_csv_dumper_1579;
    df_fifo_monitor fifo_monitor_1579;
    df_fifo_intf fifo_intf_1580(clock,reset);
    assign fifo_intf_1580.rd_en = AESL_inst_myproject.layer3_out_227_U.if_read & AESL_inst_myproject.layer3_out_227_U.if_empty_n;
    assign fifo_intf_1580.wr_en = AESL_inst_myproject.layer3_out_227_U.if_write & AESL_inst_myproject.layer3_out_227_U.if_full_n;
    assign fifo_intf_1580.fifo_rd_block = 0;
    assign fifo_intf_1580.fifo_wr_block = 0;
    assign fifo_intf_1580.finish = finish;
    csv_file_dump fifo_csv_dumper_1580;
    csv_file_dump cstatus_csv_dumper_1580;
    df_fifo_monitor fifo_monitor_1580;
    df_fifo_intf fifo_intf_1581(clock,reset);
    assign fifo_intf_1581.rd_en = AESL_inst_myproject.layer3_out_228_U.if_read & AESL_inst_myproject.layer3_out_228_U.if_empty_n;
    assign fifo_intf_1581.wr_en = AESL_inst_myproject.layer3_out_228_U.if_write & AESL_inst_myproject.layer3_out_228_U.if_full_n;
    assign fifo_intf_1581.fifo_rd_block = 0;
    assign fifo_intf_1581.fifo_wr_block = 0;
    assign fifo_intf_1581.finish = finish;
    csv_file_dump fifo_csv_dumper_1581;
    csv_file_dump cstatus_csv_dumper_1581;
    df_fifo_monitor fifo_monitor_1581;
    df_fifo_intf fifo_intf_1582(clock,reset);
    assign fifo_intf_1582.rd_en = AESL_inst_myproject.layer3_out_229_U.if_read & AESL_inst_myproject.layer3_out_229_U.if_empty_n;
    assign fifo_intf_1582.wr_en = AESL_inst_myproject.layer3_out_229_U.if_write & AESL_inst_myproject.layer3_out_229_U.if_full_n;
    assign fifo_intf_1582.fifo_rd_block = 0;
    assign fifo_intf_1582.fifo_wr_block = 0;
    assign fifo_intf_1582.finish = finish;
    csv_file_dump fifo_csv_dumper_1582;
    csv_file_dump cstatus_csv_dumper_1582;
    df_fifo_monitor fifo_monitor_1582;
    df_fifo_intf fifo_intf_1583(clock,reset);
    assign fifo_intf_1583.rd_en = AESL_inst_myproject.layer3_out_230_U.if_read & AESL_inst_myproject.layer3_out_230_U.if_empty_n;
    assign fifo_intf_1583.wr_en = AESL_inst_myproject.layer3_out_230_U.if_write & AESL_inst_myproject.layer3_out_230_U.if_full_n;
    assign fifo_intf_1583.fifo_rd_block = 0;
    assign fifo_intf_1583.fifo_wr_block = 0;
    assign fifo_intf_1583.finish = finish;
    csv_file_dump fifo_csv_dumper_1583;
    csv_file_dump cstatus_csv_dumper_1583;
    df_fifo_monitor fifo_monitor_1583;
    df_fifo_intf fifo_intf_1584(clock,reset);
    assign fifo_intf_1584.rd_en = AESL_inst_myproject.layer3_out_231_U.if_read & AESL_inst_myproject.layer3_out_231_U.if_empty_n;
    assign fifo_intf_1584.wr_en = AESL_inst_myproject.layer3_out_231_U.if_write & AESL_inst_myproject.layer3_out_231_U.if_full_n;
    assign fifo_intf_1584.fifo_rd_block = 0;
    assign fifo_intf_1584.fifo_wr_block = 0;
    assign fifo_intf_1584.finish = finish;
    csv_file_dump fifo_csv_dumper_1584;
    csv_file_dump cstatus_csv_dumper_1584;
    df_fifo_monitor fifo_monitor_1584;
    df_fifo_intf fifo_intf_1585(clock,reset);
    assign fifo_intf_1585.rd_en = AESL_inst_myproject.layer3_out_232_U.if_read & AESL_inst_myproject.layer3_out_232_U.if_empty_n;
    assign fifo_intf_1585.wr_en = AESL_inst_myproject.layer3_out_232_U.if_write & AESL_inst_myproject.layer3_out_232_U.if_full_n;
    assign fifo_intf_1585.fifo_rd_block = 0;
    assign fifo_intf_1585.fifo_wr_block = 0;
    assign fifo_intf_1585.finish = finish;
    csv_file_dump fifo_csv_dumper_1585;
    csv_file_dump cstatus_csv_dumper_1585;
    df_fifo_monitor fifo_monitor_1585;
    df_fifo_intf fifo_intf_1586(clock,reset);
    assign fifo_intf_1586.rd_en = AESL_inst_myproject.layer3_out_233_U.if_read & AESL_inst_myproject.layer3_out_233_U.if_empty_n;
    assign fifo_intf_1586.wr_en = AESL_inst_myproject.layer3_out_233_U.if_write & AESL_inst_myproject.layer3_out_233_U.if_full_n;
    assign fifo_intf_1586.fifo_rd_block = 0;
    assign fifo_intf_1586.fifo_wr_block = 0;
    assign fifo_intf_1586.finish = finish;
    csv_file_dump fifo_csv_dumper_1586;
    csv_file_dump cstatus_csv_dumper_1586;
    df_fifo_monitor fifo_monitor_1586;
    df_fifo_intf fifo_intf_1587(clock,reset);
    assign fifo_intf_1587.rd_en = AESL_inst_myproject.layer3_out_234_U.if_read & AESL_inst_myproject.layer3_out_234_U.if_empty_n;
    assign fifo_intf_1587.wr_en = AESL_inst_myproject.layer3_out_234_U.if_write & AESL_inst_myproject.layer3_out_234_U.if_full_n;
    assign fifo_intf_1587.fifo_rd_block = 0;
    assign fifo_intf_1587.fifo_wr_block = 0;
    assign fifo_intf_1587.finish = finish;
    csv_file_dump fifo_csv_dumper_1587;
    csv_file_dump cstatus_csv_dumper_1587;
    df_fifo_monitor fifo_monitor_1587;
    df_fifo_intf fifo_intf_1588(clock,reset);
    assign fifo_intf_1588.rd_en = AESL_inst_myproject.layer3_out_235_U.if_read & AESL_inst_myproject.layer3_out_235_U.if_empty_n;
    assign fifo_intf_1588.wr_en = AESL_inst_myproject.layer3_out_235_U.if_write & AESL_inst_myproject.layer3_out_235_U.if_full_n;
    assign fifo_intf_1588.fifo_rd_block = 0;
    assign fifo_intf_1588.fifo_wr_block = 0;
    assign fifo_intf_1588.finish = finish;
    csv_file_dump fifo_csv_dumper_1588;
    csv_file_dump cstatus_csv_dumper_1588;
    df_fifo_monitor fifo_monitor_1588;
    df_fifo_intf fifo_intf_1589(clock,reset);
    assign fifo_intf_1589.rd_en = AESL_inst_myproject.layer3_out_236_U.if_read & AESL_inst_myproject.layer3_out_236_U.if_empty_n;
    assign fifo_intf_1589.wr_en = AESL_inst_myproject.layer3_out_236_U.if_write & AESL_inst_myproject.layer3_out_236_U.if_full_n;
    assign fifo_intf_1589.fifo_rd_block = 0;
    assign fifo_intf_1589.fifo_wr_block = 0;
    assign fifo_intf_1589.finish = finish;
    csv_file_dump fifo_csv_dumper_1589;
    csv_file_dump cstatus_csv_dumper_1589;
    df_fifo_monitor fifo_monitor_1589;
    df_fifo_intf fifo_intf_1590(clock,reset);
    assign fifo_intf_1590.rd_en = AESL_inst_myproject.layer3_out_237_U.if_read & AESL_inst_myproject.layer3_out_237_U.if_empty_n;
    assign fifo_intf_1590.wr_en = AESL_inst_myproject.layer3_out_237_U.if_write & AESL_inst_myproject.layer3_out_237_U.if_full_n;
    assign fifo_intf_1590.fifo_rd_block = 0;
    assign fifo_intf_1590.fifo_wr_block = 0;
    assign fifo_intf_1590.finish = finish;
    csv_file_dump fifo_csv_dumper_1590;
    csv_file_dump cstatus_csv_dumper_1590;
    df_fifo_monitor fifo_monitor_1590;
    df_fifo_intf fifo_intf_1591(clock,reset);
    assign fifo_intf_1591.rd_en = AESL_inst_myproject.layer3_out_238_U.if_read & AESL_inst_myproject.layer3_out_238_U.if_empty_n;
    assign fifo_intf_1591.wr_en = AESL_inst_myproject.layer3_out_238_U.if_write & AESL_inst_myproject.layer3_out_238_U.if_full_n;
    assign fifo_intf_1591.fifo_rd_block = 0;
    assign fifo_intf_1591.fifo_wr_block = 0;
    assign fifo_intf_1591.finish = finish;
    csv_file_dump fifo_csv_dumper_1591;
    csv_file_dump cstatus_csv_dumper_1591;
    df_fifo_monitor fifo_monitor_1591;
    df_fifo_intf fifo_intf_1592(clock,reset);
    assign fifo_intf_1592.rd_en = AESL_inst_myproject.layer3_out_239_U.if_read & AESL_inst_myproject.layer3_out_239_U.if_empty_n;
    assign fifo_intf_1592.wr_en = AESL_inst_myproject.layer3_out_239_U.if_write & AESL_inst_myproject.layer3_out_239_U.if_full_n;
    assign fifo_intf_1592.fifo_rd_block = 0;
    assign fifo_intf_1592.fifo_wr_block = 0;
    assign fifo_intf_1592.finish = finish;
    csv_file_dump fifo_csv_dumper_1592;
    csv_file_dump cstatus_csv_dumper_1592;
    df_fifo_monitor fifo_monitor_1592;
    df_fifo_intf fifo_intf_1593(clock,reset);
    assign fifo_intf_1593.rd_en = AESL_inst_myproject.layer3_out_240_U.if_read & AESL_inst_myproject.layer3_out_240_U.if_empty_n;
    assign fifo_intf_1593.wr_en = AESL_inst_myproject.layer3_out_240_U.if_write & AESL_inst_myproject.layer3_out_240_U.if_full_n;
    assign fifo_intf_1593.fifo_rd_block = 0;
    assign fifo_intf_1593.fifo_wr_block = 0;
    assign fifo_intf_1593.finish = finish;
    csv_file_dump fifo_csv_dumper_1593;
    csv_file_dump cstatus_csv_dumper_1593;
    df_fifo_monitor fifo_monitor_1593;
    df_fifo_intf fifo_intf_1594(clock,reset);
    assign fifo_intf_1594.rd_en = AESL_inst_myproject.layer3_out_241_U.if_read & AESL_inst_myproject.layer3_out_241_U.if_empty_n;
    assign fifo_intf_1594.wr_en = AESL_inst_myproject.layer3_out_241_U.if_write & AESL_inst_myproject.layer3_out_241_U.if_full_n;
    assign fifo_intf_1594.fifo_rd_block = 0;
    assign fifo_intf_1594.fifo_wr_block = 0;
    assign fifo_intf_1594.finish = finish;
    csv_file_dump fifo_csv_dumper_1594;
    csv_file_dump cstatus_csv_dumper_1594;
    df_fifo_monitor fifo_monitor_1594;
    df_fifo_intf fifo_intf_1595(clock,reset);
    assign fifo_intf_1595.rd_en = AESL_inst_myproject.layer3_out_242_U.if_read & AESL_inst_myproject.layer3_out_242_U.if_empty_n;
    assign fifo_intf_1595.wr_en = AESL_inst_myproject.layer3_out_242_U.if_write & AESL_inst_myproject.layer3_out_242_U.if_full_n;
    assign fifo_intf_1595.fifo_rd_block = 0;
    assign fifo_intf_1595.fifo_wr_block = 0;
    assign fifo_intf_1595.finish = finish;
    csv_file_dump fifo_csv_dumper_1595;
    csv_file_dump cstatus_csv_dumper_1595;
    df_fifo_monitor fifo_monitor_1595;
    df_fifo_intf fifo_intf_1596(clock,reset);
    assign fifo_intf_1596.rd_en = AESL_inst_myproject.layer3_out_243_U.if_read & AESL_inst_myproject.layer3_out_243_U.if_empty_n;
    assign fifo_intf_1596.wr_en = AESL_inst_myproject.layer3_out_243_U.if_write & AESL_inst_myproject.layer3_out_243_U.if_full_n;
    assign fifo_intf_1596.fifo_rd_block = 0;
    assign fifo_intf_1596.fifo_wr_block = 0;
    assign fifo_intf_1596.finish = finish;
    csv_file_dump fifo_csv_dumper_1596;
    csv_file_dump cstatus_csv_dumper_1596;
    df_fifo_monitor fifo_monitor_1596;
    df_fifo_intf fifo_intf_1597(clock,reset);
    assign fifo_intf_1597.rd_en = AESL_inst_myproject.layer3_out_244_U.if_read & AESL_inst_myproject.layer3_out_244_U.if_empty_n;
    assign fifo_intf_1597.wr_en = AESL_inst_myproject.layer3_out_244_U.if_write & AESL_inst_myproject.layer3_out_244_U.if_full_n;
    assign fifo_intf_1597.fifo_rd_block = 0;
    assign fifo_intf_1597.fifo_wr_block = 0;
    assign fifo_intf_1597.finish = finish;
    csv_file_dump fifo_csv_dumper_1597;
    csv_file_dump cstatus_csv_dumper_1597;
    df_fifo_monitor fifo_monitor_1597;
    df_fifo_intf fifo_intf_1598(clock,reset);
    assign fifo_intf_1598.rd_en = AESL_inst_myproject.layer3_out_245_U.if_read & AESL_inst_myproject.layer3_out_245_U.if_empty_n;
    assign fifo_intf_1598.wr_en = AESL_inst_myproject.layer3_out_245_U.if_write & AESL_inst_myproject.layer3_out_245_U.if_full_n;
    assign fifo_intf_1598.fifo_rd_block = 0;
    assign fifo_intf_1598.fifo_wr_block = 0;
    assign fifo_intf_1598.finish = finish;
    csv_file_dump fifo_csv_dumper_1598;
    csv_file_dump cstatus_csv_dumper_1598;
    df_fifo_monitor fifo_monitor_1598;
    df_fifo_intf fifo_intf_1599(clock,reset);
    assign fifo_intf_1599.rd_en = AESL_inst_myproject.layer3_out_246_U.if_read & AESL_inst_myproject.layer3_out_246_U.if_empty_n;
    assign fifo_intf_1599.wr_en = AESL_inst_myproject.layer3_out_246_U.if_write & AESL_inst_myproject.layer3_out_246_U.if_full_n;
    assign fifo_intf_1599.fifo_rd_block = 0;
    assign fifo_intf_1599.fifo_wr_block = 0;
    assign fifo_intf_1599.finish = finish;
    csv_file_dump fifo_csv_dumper_1599;
    csv_file_dump cstatus_csv_dumper_1599;
    df_fifo_monitor fifo_monitor_1599;
    df_fifo_intf fifo_intf_1600(clock,reset);
    assign fifo_intf_1600.rd_en = AESL_inst_myproject.layer3_out_247_U.if_read & AESL_inst_myproject.layer3_out_247_U.if_empty_n;
    assign fifo_intf_1600.wr_en = AESL_inst_myproject.layer3_out_247_U.if_write & AESL_inst_myproject.layer3_out_247_U.if_full_n;
    assign fifo_intf_1600.fifo_rd_block = 0;
    assign fifo_intf_1600.fifo_wr_block = 0;
    assign fifo_intf_1600.finish = finish;
    csv_file_dump fifo_csv_dumper_1600;
    csv_file_dump cstatus_csv_dumper_1600;
    df_fifo_monitor fifo_monitor_1600;
    df_fifo_intf fifo_intf_1601(clock,reset);
    assign fifo_intf_1601.rd_en = AESL_inst_myproject.layer3_out_248_U.if_read & AESL_inst_myproject.layer3_out_248_U.if_empty_n;
    assign fifo_intf_1601.wr_en = AESL_inst_myproject.layer3_out_248_U.if_write & AESL_inst_myproject.layer3_out_248_U.if_full_n;
    assign fifo_intf_1601.fifo_rd_block = 0;
    assign fifo_intf_1601.fifo_wr_block = 0;
    assign fifo_intf_1601.finish = finish;
    csv_file_dump fifo_csv_dumper_1601;
    csv_file_dump cstatus_csv_dumper_1601;
    df_fifo_monitor fifo_monitor_1601;
    df_fifo_intf fifo_intf_1602(clock,reset);
    assign fifo_intf_1602.rd_en = AESL_inst_myproject.layer3_out_249_U.if_read & AESL_inst_myproject.layer3_out_249_U.if_empty_n;
    assign fifo_intf_1602.wr_en = AESL_inst_myproject.layer3_out_249_U.if_write & AESL_inst_myproject.layer3_out_249_U.if_full_n;
    assign fifo_intf_1602.fifo_rd_block = 0;
    assign fifo_intf_1602.fifo_wr_block = 0;
    assign fifo_intf_1602.finish = finish;
    csv_file_dump fifo_csv_dumper_1602;
    csv_file_dump cstatus_csv_dumper_1602;
    df_fifo_monitor fifo_monitor_1602;
    df_fifo_intf fifo_intf_1603(clock,reset);
    assign fifo_intf_1603.rd_en = AESL_inst_myproject.layer3_out_250_U.if_read & AESL_inst_myproject.layer3_out_250_U.if_empty_n;
    assign fifo_intf_1603.wr_en = AESL_inst_myproject.layer3_out_250_U.if_write & AESL_inst_myproject.layer3_out_250_U.if_full_n;
    assign fifo_intf_1603.fifo_rd_block = 0;
    assign fifo_intf_1603.fifo_wr_block = 0;
    assign fifo_intf_1603.finish = finish;
    csv_file_dump fifo_csv_dumper_1603;
    csv_file_dump cstatus_csv_dumper_1603;
    df_fifo_monitor fifo_monitor_1603;
    df_fifo_intf fifo_intf_1604(clock,reset);
    assign fifo_intf_1604.rd_en = AESL_inst_myproject.layer3_out_251_U.if_read & AESL_inst_myproject.layer3_out_251_U.if_empty_n;
    assign fifo_intf_1604.wr_en = AESL_inst_myproject.layer3_out_251_U.if_write & AESL_inst_myproject.layer3_out_251_U.if_full_n;
    assign fifo_intf_1604.fifo_rd_block = 0;
    assign fifo_intf_1604.fifo_wr_block = 0;
    assign fifo_intf_1604.finish = finish;
    csv_file_dump fifo_csv_dumper_1604;
    csv_file_dump cstatus_csv_dumper_1604;
    df_fifo_monitor fifo_monitor_1604;
    df_fifo_intf fifo_intf_1605(clock,reset);
    assign fifo_intf_1605.rd_en = AESL_inst_myproject.layer3_out_252_U.if_read & AESL_inst_myproject.layer3_out_252_U.if_empty_n;
    assign fifo_intf_1605.wr_en = AESL_inst_myproject.layer3_out_252_U.if_write & AESL_inst_myproject.layer3_out_252_U.if_full_n;
    assign fifo_intf_1605.fifo_rd_block = 0;
    assign fifo_intf_1605.fifo_wr_block = 0;
    assign fifo_intf_1605.finish = finish;
    csv_file_dump fifo_csv_dumper_1605;
    csv_file_dump cstatus_csv_dumper_1605;
    df_fifo_monitor fifo_monitor_1605;
    df_fifo_intf fifo_intf_1606(clock,reset);
    assign fifo_intf_1606.rd_en = AESL_inst_myproject.layer3_out_253_U.if_read & AESL_inst_myproject.layer3_out_253_U.if_empty_n;
    assign fifo_intf_1606.wr_en = AESL_inst_myproject.layer3_out_253_U.if_write & AESL_inst_myproject.layer3_out_253_U.if_full_n;
    assign fifo_intf_1606.fifo_rd_block = 0;
    assign fifo_intf_1606.fifo_wr_block = 0;
    assign fifo_intf_1606.finish = finish;
    csv_file_dump fifo_csv_dumper_1606;
    csv_file_dump cstatus_csv_dumper_1606;
    df_fifo_monitor fifo_monitor_1606;
    df_fifo_intf fifo_intf_1607(clock,reset);
    assign fifo_intf_1607.rd_en = AESL_inst_myproject.layer3_out_254_U.if_read & AESL_inst_myproject.layer3_out_254_U.if_empty_n;
    assign fifo_intf_1607.wr_en = AESL_inst_myproject.layer3_out_254_U.if_write & AESL_inst_myproject.layer3_out_254_U.if_full_n;
    assign fifo_intf_1607.fifo_rd_block = 0;
    assign fifo_intf_1607.fifo_wr_block = 0;
    assign fifo_intf_1607.finish = finish;
    csv_file_dump fifo_csv_dumper_1607;
    csv_file_dump cstatus_csv_dumper_1607;
    df_fifo_monitor fifo_monitor_1607;
    df_fifo_intf fifo_intf_1608(clock,reset);
    assign fifo_intf_1608.rd_en = AESL_inst_myproject.layer3_out_255_U.if_read & AESL_inst_myproject.layer3_out_255_U.if_empty_n;
    assign fifo_intf_1608.wr_en = AESL_inst_myproject.layer3_out_255_U.if_write & AESL_inst_myproject.layer3_out_255_U.if_full_n;
    assign fifo_intf_1608.fifo_rd_block = 0;
    assign fifo_intf_1608.fifo_wr_block = 0;
    assign fifo_intf_1608.finish = finish;
    csv_file_dump fifo_csv_dumper_1608;
    csv_file_dump cstatus_csv_dumper_1608;
    df_fifo_monitor fifo_monitor_1608;
    df_fifo_intf fifo_intf_1609(clock,reset);
    assign fifo_intf_1609.rd_en = AESL_inst_myproject.layer3_out_256_U.if_read & AESL_inst_myproject.layer3_out_256_U.if_empty_n;
    assign fifo_intf_1609.wr_en = AESL_inst_myproject.layer3_out_256_U.if_write & AESL_inst_myproject.layer3_out_256_U.if_full_n;
    assign fifo_intf_1609.fifo_rd_block = 0;
    assign fifo_intf_1609.fifo_wr_block = 0;
    assign fifo_intf_1609.finish = finish;
    csv_file_dump fifo_csv_dumper_1609;
    csv_file_dump cstatus_csv_dumper_1609;
    df_fifo_monitor fifo_monitor_1609;
    df_fifo_intf fifo_intf_1610(clock,reset);
    assign fifo_intf_1610.rd_en = AESL_inst_myproject.layer3_out_257_U.if_read & AESL_inst_myproject.layer3_out_257_U.if_empty_n;
    assign fifo_intf_1610.wr_en = AESL_inst_myproject.layer3_out_257_U.if_write & AESL_inst_myproject.layer3_out_257_U.if_full_n;
    assign fifo_intf_1610.fifo_rd_block = 0;
    assign fifo_intf_1610.fifo_wr_block = 0;
    assign fifo_intf_1610.finish = finish;
    csv_file_dump fifo_csv_dumper_1610;
    csv_file_dump cstatus_csv_dumper_1610;
    df_fifo_monitor fifo_monitor_1610;
    df_fifo_intf fifo_intf_1611(clock,reset);
    assign fifo_intf_1611.rd_en = AESL_inst_myproject.layer3_out_258_U.if_read & AESL_inst_myproject.layer3_out_258_U.if_empty_n;
    assign fifo_intf_1611.wr_en = AESL_inst_myproject.layer3_out_258_U.if_write & AESL_inst_myproject.layer3_out_258_U.if_full_n;
    assign fifo_intf_1611.fifo_rd_block = 0;
    assign fifo_intf_1611.fifo_wr_block = 0;
    assign fifo_intf_1611.finish = finish;
    csv_file_dump fifo_csv_dumper_1611;
    csv_file_dump cstatus_csv_dumper_1611;
    df_fifo_monitor fifo_monitor_1611;
    df_fifo_intf fifo_intf_1612(clock,reset);
    assign fifo_intf_1612.rd_en = AESL_inst_myproject.layer3_out_259_U.if_read & AESL_inst_myproject.layer3_out_259_U.if_empty_n;
    assign fifo_intf_1612.wr_en = AESL_inst_myproject.layer3_out_259_U.if_write & AESL_inst_myproject.layer3_out_259_U.if_full_n;
    assign fifo_intf_1612.fifo_rd_block = 0;
    assign fifo_intf_1612.fifo_wr_block = 0;
    assign fifo_intf_1612.finish = finish;
    csv_file_dump fifo_csv_dumper_1612;
    csv_file_dump cstatus_csv_dumper_1612;
    df_fifo_monitor fifo_monitor_1612;
    df_fifo_intf fifo_intf_1613(clock,reset);
    assign fifo_intf_1613.rd_en = AESL_inst_myproject.layer3_out_260_U.if_read & AESL_inst_myproject.layer3_out_260_U.if_empty_n;
    assign fifo_intf_1613.wr_en = AESL_inst_myproject.layer3_out_260_U.if_write & AESL_inst_myproject.layer3_out_260_U.if_full_n;
    assign fifo_intf_1613.fifo_rd_block = 0;
    assign fifo_intf_1613.fifo_wr_block = 0;
    assign fifo_intf_1613.finish = finish;
    csv_file_dump fifo_csv_dumper_1613;
    csv_file_dump cstatus_csv_dumper_1613;
    df_fifo_monitor fifo_monitor_1613;
    df_fifo_intf fifo_intf_1614(clock,reset);
    assign fifo_intf_1614.rd_en = AESL_inst_myproject.layer3_out_261_U.if_read & AESL_inst_myproject.layer3_out_261_U.if_empty_n;
    assign fifo_intf_1614.wr_en = AESL_inst_myproject.layer3_out_261_U.if_write & AESL_inst_myproject.layer3_out_261_U.if_full_n;
    assign fifo_intf_1614.fifo_rd_block = 0;
    assign fifo_intf_1614.fifo_wr_block = 0;
    assign fifo_intf_1614.finish = finish;
    csv_file_dump fifo_csv_dumper_1614;
    csv_file_dump cstatus_csv_dumper_1614;
    df_fifo_monitor fifo_monitor_1614;
    df_fifo_intf fifo_intf_1615(clock,reset);
    assign fifo_intf_1615.rd_en = AESL_inst_myproject.layer3_out_262_U.if_read & AESL_inst_myproject.layer3_out_262_U.if_empty_n;
    assign fifo_intf_1615.wr_en = AESL_inst_myproject.layer3_out_262_U.if_write & AESL_inst_myproject.layer3_out_262_U.if_full_n;
    assign fifo_intf_1615.fifo_rd_block = 0;
    assign fifo_intf_1615.fifo_wr_block = 0;
    assign fifo_intf_1615.finish = finish;
    csv_file_dump fifo_csv_dumper_1615;
    csv_file_dump cstatus_csv_dumper_1615;
    df_fifo_monitor fifo_monitor_1615;
    df_fifo_intf fifo_intf_1616(clock,reset);
    assign fifo_intf_1616.rd_en = AESL_inst_myproject.layer3_out_263_U.if_read & AESL_inst_myproject.layer3_out_263_U.if_empty_n;
    assign fifo_intf_1616.wr_en = AESL_inst_myproject.layer3_out_263_U.if_write & AESL_inst_myproject.layer3_out_263_U.if_full_n;
    assign fifo_intf_1616.fifo_rd_block = 0;
    assign fifo_intf_1616.fifo_wr_block = 0;
    assign fifo_intf_1616.finish = finish;
    csv_file_dump fifo_csv_dumper_1616;
    csv_file_dump cstatus_csv_dumper_1616;
    df_fifo_monitor fifo_monitor_1616;
    df_fifo_intf fifo_intf_1617(clock,reset);
    assign fifo_intf_1617.rd_en = AESL_inst_myproject.layer3_out_264_U.if_read & AESL_inst_myproject.layer3_out_264_U.if_empty_n;
    assign fifo_intf_1617.wr_en = AESL_inst_myproject.layer3_out_264_U.if_write & AESL_inst_myproject.layer3_out_264_U.if_full_n;
    assign fifo_intf_1617.fifo_rd_block = 0;
    assign fifo_intf_1617.fifo_wr_block = 0;
    assign fifo_intf_1617.finish = finish;
    csv_file_dump fifo_csv_dumper_1617;
    csv_file_dump cstatus_csv_dumper_1617;
    df_fifo_monitor fifo_monitor_1617;
    df_fifo_intf fifo_intf_1618(clock,reset);
    assign fifo_intf_1618.rd_en = AESL_inst_myproject.layer3_out_265_U.if_read & AESL_inst_myproject.layer3_out_265_U.if_empty_n;
    assign fifo_intf_1618.wr_en = AESL_inst_myproject.layer3_out_265_U.if_write & AESL_inst_myproject.layer3_out_265_U.if_full_n;
    assign fifo_intf_1618.fifo_rd_block = 0;
    assign fifo_intf_1618.fifo_wr_block = 0;
    assign fifo_intf_1618.finish = finish;
    csv_file_dump fifo_csv_dumper_1618;
    csv_file_dump cstatus_csv_dumper_1618;
    df_fifo_monitor fifo_monitor_1618;
    df_fifo_intf fifo_intf_1619(clock,reset);
    assign fifo_intf_1619.rd_en = AESL_inst_myproject.layer3_out_266_U.if_read & AESL_inst_myproject.layer3_out_266_U.if_empty_n;
    assign fifo_intf_1619.wr_en = AESL_inst_myproject.layer3_out_266_U.if_write & AESL_inst_myproject.layer3_out_266_U.if_full_n;
    assign fifo_intf_1619.fifo_rd_block = 0;
    assign fifo_intf_1619.fifo_wr_block = 0;
    assign fifo_intf_1619.finish = finish;
    csv_file_dump fifo_csv_dumper_1619;
    csv_file_dump cstatus_csv_dumper_1619;
    df_fifo_monitor fifo_monitor_1619;
    df_fifo_intf fifo_intf_1620(clock,reset);
    assign fifo_intf_1620.rd_en = AESL_inst_myproject.layer3_out_267_U.if_read & AESL_inst_myproject.layer3_out_267_U.if_empty_n;
    assign fifo_intf_1620.wr_en = AESL_inst_myproject.layer3_out_267_U.if_write & AESL_inst_myproject.layer3_out_267_U.if_full_n;
    assign fifo_intf_1620.fifo_rd_block = 0;
    assign fifo_intf_1620.fifo_wr_block = 0;
    assign fifo_intf_1620.finish = finish;
    csv_file_dump fifo_csv_dumper_1620;
    csv_file_dump cstatus_csv_dumper_1620;
    df_fifo_monitor fifo_monitor_1620;
    df_fifo_intf fifo_intf_1621(clock,reset);
    assign fifo_intf_1621.rd_en = AESL_inst_myproject.layer3_out_268_U.if_read & AESL_inst_myproject.layer3_out_268_U.if_empty_n;
    assign fifo_intf_1621.wr_en = AESL_inst_myproject.layer3_out_268_U.if_write & AESL_inst_myproject.layer3_out_268_U.if_full_n;
    assign fifo_intf_1621.fifo_rd_block = 0;
    assign fifo_intf_1621.fifo_wr_block = 0;
    assign fifo_intf_1621.finish = finish;
    csv_file_dump fifo_csv_dumper_1621;
    csv_file_dump cstatus_csv_dumper_1621;
    df_fifo_monitor fifo_monitor_1621;
    df_fifo_intf fifo_intf_1622(clock,reset);
    assign fifo_intf_1622.rd_en = AESL_inst_myproject.layer3_out_269_U.if_read & AESL_inst_myproject.layer3_out_269_U.if_empty_n;
    assign fifo_intf_1622.wr_en = AESL_inst_myproject.layer3_out_269_U.if_write & AESL_inst_myproject.layer3_out_269_U.if_full_n;
    assign fifo_intf_1622.fifo_rd_block = 0;
    assign fifo_intf_1622.fifo_wr_block = 0;
    assign fifo_intf_1622.finish = finish;
    csv_file_dump fifo_csv_dumper_1622;
    csv_file_dump cstatus_csv_dumper_1622;
    df_fifo_monitor fifo_monitor_1622;
    df_fifo_intf fifo_intf_1623(clock,reset);
    assign fifo_intf_1623.rd_en = AESL_inst_myproject.layer3_out_270_U.if_read & AESL_inst_myproject.layer3_out_270_U.if_empty_n;
    assign fifo_intf_1623.wr_en = AESL_inst_myproject.layer3_out_270_U.if_write & AESL_inst_myproject.layer3_out_270_U.if_full_n;
    assign fifo_intf_1623.fifo_rd_block = 0;
    assign fifo_intf_1623.fifo_wr_block = 0;
    assign fifo_intf_1623.finish = finish;
    csv_file_dump fifo_csv_dumper_1623;
    csv_file_dump cstatus_csv_dumper_1623;
    df_fifo_monitor fifo_monitor_1623;
    df_fifo_intf fifo_intf_1624(clock,reset);
    assign fifo_intf_1624.rd_en = AESL_inst_myproject.layer3_out_271_U.if_read & AESL_inst_myproject.layer3_out_271_U.if_empty_n;
    assign fifo_intf_1624.wr_en = AESL_inst_myproject.layer3_out_271_U.if_write & AESL_inst_myproject.layer3_out_271_U.if_full_n;
    assign fifo_intf_1624.fifo_rd_block = 0;
    assign fifo_intf_1624.fifo_wr_block = 0;
    assign fifo_intf_1624.finish = finish;
    csv_file_dump fifo_csv_dumper_1624;
    csv_file_dump cstatus_csv_dumper_1624;
    df_fifo_monitor fifo_monitor_1624;
    df_fifo_intf fifo_intf_1625(clock,reset);
    assign fifo_intf_1625.rd_en = AESL_inst_myproject.layer3_out_272_U.if_read & AESL_inst_myproject.layer3_out_272_U.if_empty_n;
    assign fifo_intf_1625.wr_en = AESL_inst_myproject.layer3_out_272_U.if_write & AESL_inst_myproject.layer3_out_272_U.if_full_n;
    assign fifo_intf_1625.fifo_rd_block = 0;
    assign fifo_intf_1625.fifo_wr_block = 0;
    assign fifo_intf_1625.finish = finish;
    csv_file_dump fifo_csv_dumper_1625;
    csv_file_dump cstatus_csv_dumper_1625;
    df_fifo_monitor fifo_monitor_1625;
    df_fifo_intf fifo_intf_1626(clock,reset);
    assign fifo_intf_1626.rd_en = AESL_inst_myproject.layer3_out_273_U.if_read & AESL_inst_myproject.layer3_out_273_U.if_empty_n;
    assign fifo_intf_1626.wr_en = AESL_inst_myproject.layer3_out_273_U.if_write & AESL_inst_myproject.layer3_out_273_U.if_full_n;
    assign fifo_intf_1626.fifo_rd_block = 0;
    assign fifo_intf_1626.fifo_wr_block = 0;
    assign fifo_intf_1626.finish = finish;
    csv_file_dump fifo_csv_dumper_1626;
    csv_file_dump cstatus_csv_dumper_1626;
    df_fifo_monitor fifo_monitor_1626;
    df_fifo_intf fifo_intf_1627(clock,reset);
    assign fifo_intf_1627.rd_en = AESL_inst_myproject.layer3_out_274_U.if_read & AESL_inst_myproject.layer3_out_274_U.if_empty_n;
    assign fifo_intf_1627.wr_en = AESL_inst_myproject.layer3_out_274_U.if_write & AESL_inst_myproject.layer3_out_274_U.if_full_n;
    assign fifo_intf_1627.fifo_rd_block = 0;
    assign fifo_intf_1627.fifo_wr_block = 0;
    assign fifo_intf_1627.finish = finish;
    csv_file_dump fifo_csv_dumper_1627;
    csv_file_dump cstatus_csv_dumper_1627;
    df_fifo_monitor fifo_monitor_1627;
    df_fifo_intf fifo_intf_1628(clock,reset);
    assign fifo_intf_1628.rd_en = AESL_inst_myproject.layer3_out_275_U.if_read & AESL_inst_myproject.layer3_out_275_U.if_empty_n;
    assign fifo_intf_1628.wr_en = AESL_inst_myproject.layer3_out_275_U.if_write & AESL_inst_myproject.layer3_out_275_U.if_full_n;
    assign fifo_intf_1628.fifo_rd_block = 0;
    assign fifo_intf_1628.fifo_wr_block = 0;
    assign fifo_intf_1628.finish = finish;
    csv_file_dump fifo_csv_dumper_1628;
    csv_file_dump cstatus_csv_dumper_1628;
    df_fifo_monitor fifo_monitor_1628;
    df_fifo_intf fifo_intf_1629(clock,reset);
    assign fifo_intf_1629.rd_en = AESL_inst_myproject.layer3_out_276_U.if_read & AESL_inst_myproject.layer3_out_276_U.if_empty_n;
    assign fifo_intf_1629.wr_en = AESL_inst_myproject.layer3_out_276_U.if_write & AESL_inst_myproject.layer3_out_276_U.if_full_n;
    assign fifo_intf_1629.fifo_rd_block = 0;
    assign fifo_intf_1629.fifo_wr_block = 0;
    assign fifo_intf_1629.finish = finish;
    csv_file_dump fifo_csv_dumper_1629;
    csv_file_dump cstatus_csv_dumper_1629;
    df_fifo_monitor fifo_monitor_1629;
    df_fifo_intf fifo_intf_1630(clock,reset);
    assign fifo_intf_1630.rd_en = AESL_inst_myproject.layer3_out_277_U.if_read & AESL_inst_myproject.layer3_out_277_U.if_empty_n;
    assign fifo_intf_1630.wr_en = AESL_inst_myproject.layer3_out_277_U.if_write & AESL_inst_myproject.layer3_out_277_U.if_full_n;
    assign fifo_intf_1630.fifo_rd_block = 0;
    assign fifo_intf_1630.fifo_wr_block = 0;
    assign fifo_intf_1630.finish = finish;
    csv_file_dump fifo_csv_dumper_1630;
    csv_file_dump cstatus_csv_dumper_1630;
    df_fifo_monitor fifo_monitor_1630;
    df_fifo_intf fifo_intf_1631(clock,reset);
    assign fifo_intf_1631.rd_en = AESL_inst_myproject.layer3_out_278_U.if_read & AESL_inst_myproject.layer3_out_278_U.if_empty_n;
    assign fifo_intf_1631.wr_en = AESL_inst_myproject.layer3_out_278_U.if_write & AESL_inst_myproject.layer3_out_278_U.if_full_n;
    assign fifo_intf_1631.fifo_rd_block = 0;
    assign fifo_intf_1631.fifo_wr_block = 0;
    assign fifo_intf_1631.finish = finish;
    csv_file_dump fifo_csv_dumper_1631;
    csv_file_dump cstatus_csv_dumper_1631;
    df_fifo_monitor fifo_monitor_1631;
    df_fifo_intf fifo_intf_1632(clock,reset);
    assign fifo_intf_1632.rd_en = AESL_inst_myproject.layer3_out_279_U.if_read & AESL_inst_myproject.layer3_out_279_U.if_empty_n;
    assign fifo_intf_1632.wr_en = AESL_inst_myproject.layer3_out_279_U.if_write & AESL_inst_myproject.layer3_out_279_U.if_full_n;
    assign fifo_intf_1632.fifo_rd_block = 0;
    assign fifo_intf_1632.fifo_wr_block = 0;
    assign fifo_intf_1632.finish = finish;
    csv_file_dump fifo_csv_dumper_1632;
    csv_file_dump cstatus_csv_dumper_1632;
    df_fifo_monitor fifo_monitor_1632;
    df_fifo_intf fifo_intf_1633(clock,reset);
    assign fifo_intf_1633.rd_en = AESL_inst_myproject.layer3_out_280_U.if_read & AESL_inst_myproject.layer3_out_280_U.if_empty_n;
    assign fifo_intf_1633.wr_en = AESL_inst_myproject.layer3_out_280_U.if_write & AESL_inst_myproject.layer3_out_280_U.if_full_n;
    assign fifo_intf_1633.fifo_rd_block = 0;
    assign fifo_intf_1633.fifo_wr_block = 0;
    assign fifo_intf_1633.finish = finish;
    csv_file_dump fifo_csv_dumper_1633;
    csv_file_dump cstatus_csv_dumper_1633;
    df_fifo_monitor fifo_monitor_1633;
    df_fifo_intf fifo_intf_1634(clock,reset);
    assign fifo_intf_1634.rd_en = AESL_inst_myproject.layer3_out_281_U.if_read & AESL_inst_myproject.layer3_out_281_U.if_empty_n;
    assign fifo_intf_1634.wr_en = AESL_inst_myproject.layer3_out_281_U.if_write & AESL_inst_myproject.layer3_out_281_U.if_full_n;
    assign fifo_intf_1634.fifo_rd_block = 0;
    assign fifo_intf_1634.fifo_wr_block = 0;
    assign fifo_intf_1634.finish = finish;
    csv_file_dump fifo_csv_dumper_1634;
    csv_file_dump cstatus_csv_dumper_1634;
    df_fifo_monitor fifo_monitor_1634;
    df_fifo_intf fifo_intf_1635(clock,reset);
    assign fifo_intf_1635.rd_en = AESL_inst_myproject.layer3_out_282_U.if_read & AESL_inst_myproject.layer3_out_282_U.if_empty_n;
    assign fifo_intf_1635.wr_en = AESL_inst_myproject.layer3_out_282_U.if_write & AESL_inst_myproject.layer3_out_282_U.if_full_n;
    assign fifo_intf_1635.fifo_rd_block = 0;
    assign fifo_intf_1635.fifo_wr_block = 0;
    assign fifo_intf_1635.finish = finish;
    csv_file_dump fifo_csv_dumper_1635;
    csv_file_dump cstatus_csv_dumper_1635;
    df_fifo_monitor fifo_monitor_1635;
    df_fifo_intf fifo_intf_1636(clock,reset);
    assign fifo_intf_1636.rd_en = AESL_inst_myproject.layer3_out_283_U.if_read & AESL_inst_myproject.layer3_out_283_U.if_empty_n;
    assign fifo_intf_1636.wr_en = AESL_inst_myproject.layer3_out_283_U.if_write & AESL_inst_myproject.layer3_out_283_U.if_full_n;
    assign fifo_intf_1636.fifo_rd_block = 0;
    assign fifo_intf_1636.fifo_wr_block = 0;
    assign fifo_intf_1636.finish = finish;
    csv_file_dump fifo_csv_dumper_1636;
    csv_file_dump cstatus_csv_dumper_1636;
    df_fifo_monitor fifo_monitor_1636;
    df_fifo_intf fifo_intf_1637(clock,reset);
    assign fifo_intf_1637.rd_en = AESL_inst_myproject.layer3_out_284_U.if_read & AESL_inst_myproject.layer3_out_284_U.if_empty_n;
    assign fifo_intf_1637.wr_en = AESL_inst_myproject.layer3_out_284_U.if_write & AESL_inst_myproject.layer3_out_284_U.if_full_n;
    assign fifo_intf_1637.fifo_rd_block = 0;
    assign fifo_intf_1637.fifo_wr_block = 0;
    assign fifo_intf_1637.finish = finish;
    csv_file_dump fifo_csv_dumper_1637;
    csv_file_dump cstatus_csv_dumper_1637;
    df_fifo_monitor fifo_monitor_1637;
    df_fifo_intf fifo_intf_1638(clock,reset);
    assign fifo_intf_1638.rd_en = AESL_inst_myproject.layer3_out_285_U.if_read & AESL_inst_myproject.layer3_out_285_U.if_empty_n;
    assign fifo_intf_1638.wr_en = AESL_inst_myproject.layer3_out_285_U.if_write & AESL_inst_myproject.layer3_out_285_U.if_full_n;
    assign fifo_intf_1638.fifo_rd_block = 0;
    assign fifo_intf_1638.fifo_wr_block = 0;
    assign fifo_intf_1638.finish = finish;
    csv_file_dump fifo_csv_dumper_1638;
    csv_file_dump cstatus_csv_dumper_1638;
    df_fifo_monitor fifo_monitor_1638;
    df_fifo_intf fifo_intf_1639(clock,reset);
    assign fifo_intf_1639.rd_en = AESL_inst_myproject.layer3_out_286_U.if_read & AESL_inst_myproject.layer3_out_286_U.if_empty_n;
    assign fifo_intf_1639.wr_en = AESL_inst_myproject.layer3_out_286_U.if_write & AESL_inst_myproject.layer3_out_286_U.if_full_n;
    assign fifo_intf_1639.fifo_rd_block = 0;
    assign fifo_intf_1639.fifo_wr_block = 0;
    assign fifo_intf_1639.finish = finish;
    csv_file_dump fifo_csv_dumper_1639;
    csv_file_dump cstatus_csv_dumper_1639;
    df_fifo_monitor fifo_monitor_1639;
    df_fifo_intf fifo_intf_1640(clock,reset);
    assign fifo_intf_1640.rd_en = AESL_inst_myproject.layer3_out_287_U.if_read & AESL_inst_myproject.layer3_out_287_U.if_empty_n;
    assign fifo_intf_1640.wr_en = AESL_inst_myproject.layer3_out_287_U.if_write & AESL_inst_myproject.layer3_out_287_U.if_full_n;
    assign fifo_intf_1640.fifo_rd_block = 0;
    assign fifo_intf_1640.fifo_wr_block = 0;
    assign fifo_intf_1640.finish = finish;
    csv_file_dump fifo_csv_dumper_1640;
    csv_file_dump cstatus_csv_dumper_1640;
    df_fifo_monitor fifo_monitor_1640;
    df_fifo_intf fifo_intf_1641(clock,reset);
    assign fifo_intf_1641.rd_en = AESL_inst_myproject.layer3_out_288_U.if_read & AESL_inst_myproject.layer3_out_288_U.if_empty_n;
    assign fifo_intf_1641.wr_en = AESL_inst_myproject.layer3_out_288_U.if_write & AESL_inst_myproject.layer3_out_288_U.if_full_n;
    assign fifo_intf_1641.fifo_rd_block = 0;
    assign fifo_intf_1641.fifo_wr_block = 0;
    assign fifo_intf_1641.finish = finish;
    csv_file_dump fifo_csv_dumper_1641;
    csv_file_dump cstatus_csv_dumper_1641;
    df_fifo_monitor fifo_monitor_1641;
    df_fifo_intf fifo_intf_1642(clock,reset);
    assign fifo_intf_1642.rd_en = AESL_inst_myproject.layer3_out_289_U.if_read & AESL_inst_myproject.layer3_out_289_U.if_empty_n;
    assign fifo_intf_1642.wr_en = AESL_inst_myproject.layer3_out_289_U.if_write & AESL_inst_myproject.layer3_out_289_U.if_full_n;
    assign fifo_intf_1642.fifo_rd_block = 0;
    assign fifo_intf_1642.fifo_wr_block = 0;
    assign fifo_intf_1642.finish = finish;
    csv_file_dump fifo_csv_dumper_1642;
    csv_file_dump cstatus_csv_dumper_1642;
    df_fifo_monitor fifo_monitor_1642;
    df_fifo_intf fifo_intf_1643(clock,reset);
    assign fifo_intf_1643.rd_en = AESL_inst_myproject.layer3_out_290_U.if_read & AESL_inst_myproject.layer3_out_290_U.if_empty_n;
    assign fifo_intf_1643.wr_en = AESL_inst_myproject.layer3_out_290_U.if_write & AESL_inst_myproject.layer3_out_290_U.if_full_n;
    assign fifo_intf_1643.fifo_rd_block = 0;
    assign fifo_intf_1643.fifo_wr_block = 0;
    assign fifo_intf_1643.finish = finish;
    csv_file_dump fifo_csv_dumper_1643;
    csv_file_dump cstatus_csv_dumper_1643;
    df_fifo_monitor fifo_monitor_1643;
    df_fifo_intf fifo_intf_1644(clock,reset);
    assign fifo_intf_1644.rd_en = AESL_inst_myproject.layer3_out_291_U.if_read & AESL_inst_myproject.layer3_out_291_U.if_empty_n;
    assign fifo_intf_1644.wr_en = AESL_inst_myproject.layer3_out_291_U.if_write & AESL_inst_myproject.layer3_out_291_U.if_full_n;
    assign fifo_intf_1644.fifo_rd_block = 0;
    assign fifo_intf_1644.fifo_wr_block = 0;
    assign fifo_intf_1644.finish = finish;
    csv_file_dump fifo_csv_dumper_1644;
    csv_file_dump cstatus_csv_dumper_1644;
    df_fifo_monitor fifo_monitor_1644;
    df_fifo_intf fifo_intf_1645(clock,reset);
    assign fifo_intf_1645.rd_en = AESL_inst_myproject.layer3_out_292_U.if_read & AESL_inst_myproject.layer3_out_292_U.if_empty_n;
    assign fifo_intf_1645.wr_en = AESL_inst_myproject.layer3_out_292_U.if_write & AESL_inst_myproject.layer3_out_292_U.if_full_n;
    assign fifo_intf_1645.fifo_rd_block = 0;
    assign fifo_intf_1645.fifo_wr_block = 0;
    assign fifo_intf_1645.finish = finish;
    csv_file_dump fifo_csv_dumper_1645;
    csv_file_dump cstatus_csv_dumper_1645;
    df_fifo_monitor fifo_monitor_1645;
    df_fifo_intf fifo_intf_1646(clock,reset);
    assign fifo_intf_1646.rd_en = AESL_inst_myproject.layer3_out_293_U.if_read & AESL_inst_myproject.layer3_out_293_U.if_empty_n;
    assign fifo_intf_1646.wr_en = AESL_inst_myproject.layer3_out_293_U.if_write & AESL_inst_myproject.layer3_out_293_U.if_full_n;
    assign fifo_intf_1646.fifo_rd_block = 0;
    assign fifo_intf_1646.fifo_wr_block = 0;
    assign fifo_intf_1646.finish = finish;
    csv_file_dump fifo_csv_dumper_1646;
    csv_file_dump cstatus_csv_dumper_1646;
    df_fifo_monitor fifo_monitor_1646;
    df_fifo_intf fifo_intf_1647(clock,reset);
    assign fifo_intf_1647.rd_en = AESL_inst_myproject.layer3_out_294_U.if_read & AESL_inst_myproject.layer3_out_294_U.if_empty_n;
    assign fifo_intf_1647.wr_en = AESL_inst_myproject.layer3_out_294_U.if_write & AESL_inst_myproject.layer3_out_294_U.if_full_n;
    assign fifo_intf_1647.fifo_rd_block = 0;
    assign fifo_intf_1647.fifo_wr_block = 0;
    assign fifo_intf_1647.finish = finish;
    csv_file_dump fifo_csv_dumper_1647;
    csv_file_dump cstatus_csv_dumper_1647;
    df_fifo_monitor fifo_monitor_1647;
    df_fifo_intf fifo_intf_1648(clock,reset);
    assign fifo_intf_1648.rd_en = AESL_inst_myproject.layer3_out_295_U.if_read & AESL_inst_myproject.layer3_out_295_U.if_empty_n;
    assign fifo_intf_1648.wr_en = AESL_inst_myproject.layer3_out_295_U.if_write & AESL_inst_myproject.layer3_out_295_U.if_full_n;
    assign fifo_intf_1648.fifo_rd_block = 0;
    assign fifo_intf_1648.fifo_wr_block = 0;
    assign fifo_intf_1648.finish = finish;
    csv_file_dump fifo_csv_dumper_1648;
    csv_file_dump cstatus_csv_dumper_1648;
    df_fifo_monitor fifo_monitor_1648;
    df_fifo_intf fifo_intf_1649(clock,reset);
    assign fifo_intf_1649.rd_en = AESL_inst_myproject.layer3_out_296_U.if_read & AESL_inst_myproject.layer3_out_296_U.if_empty_n;
    assign fifo_intf_1649.wr_en = AESL_inst_myproject.layer3_out_296_U.if_write & AESL_inst_myproject.layer3_out_296_U.if_full_n;
    assign fifo_intf_1649.fifo_rd_block = 0;
    assign fifo_intf_1649.fifo_wr_block = 0;
    assign fifo_intf_1649.finish = finish;
    csv_file_dump fifo_csv_dumper_1649;
    csv_file_dump cstatus_csv_dumper_1649;
    df_fifo_monitor fifo_monitor_1649;
    df_fifo_intf fifo_intf_1650(clock,reset);
    assign fifo_intf_1650.rd_en = AESL_inst_myproject.layer3_out_297_U.if_read & AESL_inst_myproject.layer3_out_297_U.if_empty_n;
    assign fifo_intf_1650.wr_en = AESL_inst_myproject.layer3_out_297_U.if_write & AESL_inst_myproject.layer3_out_297_U.if_full_n;
    assign fifo_intf_1650.fifo_rd_block = 0;
    assign fifo_intf_1650.fifo_wr_block = 0;
    assign fifo_intf_1650.finish = finish;
    csv_file_dump fifo_csv_dumper_1650;
    csv_file_dump cstatus_csv_dumper_1650;
    df_fifo_monitor fifo_monitor_1650;
    df_fifo_intf fifo_intf_1651(clock,reset);
    assign fifo_intf_1651.rd_en = AESL_inst_myproject.layer3_out_298_U.if_read & AESL_inst_myproject.layer3_out_298_U.if_empty_n;
    assign fifo_intf_1651.wr_en = AESL_inst_myproject.layer3_out_298_U.if_write & AESL_inst_myproject.layer3_out_298_U.if_full_n;
    assign fifo_intf_1651.fifo_rd_block = 0;
    assign fifo_intf_1651.fifo_wr_block = 0;
    assign fifo_intf_1651.finish = finish;
    csv_file_dump fifo_csv_dumper_1651;
    csv_file_dump cstatus_csv_dumper_1651;
    df_fifo_monitor fifo_monitor_1651;
    df_fifo_intf fifo_intf_1652(clock,reset);
    assign fifo_intf_1652.rd_en = AESL_inst_myproject.layer3_out_299_U.if_read & AESL_inst_myproject.layer3_out_299_U.if_empty_n;
    assign fifo_intf_1652.wr_en = AESL_inst_myproject.layer3_out_299_U.if_write & AESL_inst_myproject.layer3_out_299_U.if_full_n;
    assign fifo_intf_1652.fifo_rd_block = 0;
    assign fifo_intf_1652.fifo_wr_block = 0;
    assign fifo_intf_1652.finish = finish;
    csv_file_dump fifo_csv_dumper_1652;
    csv_file_dump cstatus_csv_dumper_1652;
    df_fifo_monitor fifo_monitor_1652;
    df_fifo_intf fifo_intf_1653(clock,reset);
    assign fifo_intf_1653.rd_en = AESL_inst_myproject.layer3_out_300_U.if_read & AESL_inst_myproject.layer3_out_300_U.if_empty_n;
    assign fifo_intf_1653.wr_en = AESL_inst_myproject.layer3_out_300_U.if_write & AESL_inst_myproject.layer3_out_300_U.if_full_n;
    assign fifo_intf_1653.fifo_rd_block = 0;
    assign fifo_intf_1653.fifo_wr_block = 0;
    assign fifo_intf_1653.finish = finish;
    csv_file_dump fifo_csv_dumper_1653;
    csv_file_dump cstatus_csv_dumper_1653;
    df_fifo_monitor fifo_monitor_1653;
    df_fifo_intf fifo_intf_1654(clock,reset);
    assign fifo_intf_1654.rd_en = AESL_inst_myproject.layer3_out_301_U.if_read & AESL_inst_myproject.layer3_out_301_U.if_empty_n;
    assign fifo_intf_1654.wr_en = AESL_inst_myproject.layer3_out_301_U.if_write & AESL_inst_myproject.layer3_out_301_U.if_full_n;
    assign fifo_intf_1654.fifo_rd_block = 0;
    assign fifo_intf_1654.fifo_wr_block = 0;
    assign fifo_intf_1654.finish = finish;
    csv_file_dump fifo_csv_dumper_1654;
    csv_file_dump cstatus_csv_dumper_1654;
    df_fifo_monitor fifo_monitor_1654;
    df_fifo_intf fifo_intf_1655(clock,reset);
    assign fifo_intf_1655.rd_en = AESL_inst_myproject.layer3_out_302_U.if_read & AESL_inst_myproject.layer3_out_302_U.if_empty_n;
    assign fifo_intf_1655.wr_en = AESL_inst_myproject.layer3_out_302_U.if_write & AESL_inst_myproject.layer3_out_302_U.if_full_n;
    assign fifo_intf_1655.fifo_rd_block = 0;
    assign fifo_intf_1655.fifo_wr_block = 0;
    assign fifo_intf_1655.finish = finish;
    csv_file_dump fifo_csv_dumper_1655;
    csv_file_dump cstatus_csv_dumper_1655;
    df_fifo_monitor fifo_monitor_1655;
    df_fifo_intf fifo_intf_1656(clock,reset);
    assign fifo_intf_1656.rd_en = AESL_inst_myproject.layer3_out_303_U.if_read & AESL_inst_myproject.layer3_out_303_U.if_empty_n;
    assign fifo_intf_1656.wr_en = AESL_inst_myproject.layer3_out_303_U.if_write & AESL_inst_myproject.layer3_out_303_U.if_full_n;
    assign fifo_intf_1656.fifo_rd_block = 0;
    assign fifo_intf_1656.fifo_wr_block = 0;
    assign fifo_intf_1656.finish = finish;
    csv_file_dump fifo_csv_dumper_1656;
    csv_file_dump cstatus_csv_dumper_1656;
    df_fifo_monitor fifo_monitor_1656;
    df_fifo_intf fifo_intf_1657(clock,reset);
    assign fifo_intf_1657.rd_en = AESL_inst_myproject.layer3_out_304_U.if_read & AESL_inst_myproject.layer3_out_304_U.if_empty_n;
    assign fifo_intf_1657.wr_en = AESL_inst_myproject.layer3_out_304_U.if_write & AESL_inst_myproject.layer3_out_304_U.if_full_n;
    assign fifo_intf_1657.fifo_rd_block = 0;
    assign fifo_intf_1657.fifo_wr_block = 0;
    assign fifo_intf_1657.finish = finish;
    csv_file_dump fifo_csv_dumper_1657;
    csv_file_dump cstatus_csv_dumper_1657;
    df_fifo_monitor fifo_monitor_1657;
    df_fifo_intf fifo_intf_1658(clock,reset);
    assign fifo_intf_1658.rd_en = AESL_inst_myproject.layer3_out_305_U.if_read & AESL_inst_myproject.layer3_out_305_U.if_empty_n;
    assign fifo_intf_1658.wr_en = AESL_inst_myproject.layer3_out_305_U.if_write & AESL_inst_myproject.layer3_out_305_U.if_full_n;
    assign fifo_intf_1658.fifo_rd_block = 0;
    assign fifo_intf_1658.fifo_wr_block = 0;
    assign fifo_intf_1658.finish = finish;
    csv_file_dump fifo_csv_dumper_1658;
    csv_file_dump cstatus_csv_dumper_1658;
    df_fifo_monitor fifo_monitor_1658;
    df_fifo_intf fifo_intf_1659(clock,reset);
    assign fifo_intf_1659.rd_en = AESL_inst_myproject.layer3_out_306_U.if_read & AESL_inst_myproject.layer3_out_306_U.if_empty_n;
    assign fifo_intf_1659.wr_en = AESL_inst_myproject.layer3_out_306_U.if_write & AESL_inst_myproject.layer3_out_306_U.if_full_n;
    assign fifo_intf_1659.fifo_rd_block = 0;
    assign fifo_intf_1659.fifo_wr_block = 0;
    assign fifo_intf_1659.finish = finish;
    csv_file_dump fifo_csv_dumper_1659;
    csv_file_dump cstatus_csv_dumper_1659;
    df_fifo_monitor fifo_monitor_1659;
    df_fifo_intf fifo_intf_1660(clock,reset);
    assign fifo_intf_1660.rd_en = AESL_inst_myproject.layer3_out_307_U.if_read & AESL_inst_myproject.layer3_out_307_U.if_empty_n;
    assign fifo_intf_1660.wr_en = AESL_inst_myproject.layer3_out_307_U.if_write & AESL_inst_myproject.layer3_out_307_U.if_full_n;
    assign fifo_intf_1660.fifo_rd_block = 0;
    assign fifo_intf_1660.fifo_wr_block = 0;
    assign fifo_intf_1660.finish = finish;
    csv_file_dump fifo_csv_dumper_1660;
    csv_file_dump cstatus_csv_dumper_1660;
    df_fifo_monitor fifo_monitor_1660;
    df_fifo_intf fifo_intf_1661(clock,reset);
    assign fifo_intf_1661.rd_en = AESL_inst_myproject.layer3_out_308_U.if_read & AESL_inst_myproject.layer3_out_308_U.if_empty_n;
    assign fifo_intf_1661.wr_en = AESL_inst_myproject.layer3_out_308_U.if_write & AESL_inst_myproject.layer3_out_308_U.if_full_n;
    assign fifo_intf_1661.fifo_rd_block = 0;
    assign fifo_intf_1661.fifo_wr_block = 0;
    assign fifo_intf_1661.finish = finish;
    csv_file_dump fifo_csv_dumper_1661;
    csv_file_dump cstatus_csv_dumper_1661;
    df_fifo_monitor fifo_monitor_1661;
    df_fifo_intf fifo_intf_1662(clock,reset);
    assign fifo_intf_1662.rd_en = AESL_inst_myproject.layer3_out_309_U.if_read & AESL_inst_myproject.layer3_out_309_U.if_empty_n;
    assign fifo_intf_1662.wr_en = AESL_inst_myproject.layer3_out_309_U.if_write & AESL_inst_myproject.layer3_out_309_U.if_full_n;
    assign fifo_intf_1662.fifo_rd_block = 0;
    assign fifo_intf_1662.fifo_wr_block = 0;
    assign fifo_intf_1662.finish = finish;
    csv_file_dump fifo_csv_dumper_1662;
    csv_file_dump cstatus_csv_dumper_1662;
    df_fifo_monitor fifo_monitor_1662;
    df_fifo_intf fifo_intf_1663(clock,reset);
    assign fifo_intf_1663.rd_en = AESL_inst_myproject.layer3_out_310_U.if_read & AESL_inst_myproject.layer3_out_310_U.if_empty_n;
    assign fifo_intf_1663.wr_en = AESL_inst_myproject.layer3_out_310_U.if_write & AESL_inst_myproject.layer3_out_310_U.if_full_n;
    assign fifo_intf_1663.fifo_rd_block = 0;
    assign fifo_intf_1663.fifo_wr_block = 0;
    assign fifo_intf_1663.finish = finish;
    csv_file_dump fifo_csv_dumper_1663;
    csv_file_dump cstatus_csv_dumper_1663;
    df_fifo_monitor fifo_monitor_1663;
    df_fifo_intf fifo_intf_1664(clock,reset);
    assign fifo_intf_1664.rd_en = AESL_inst_myproject.layer3_out_311_U.if_read & AESL_inst_myproject.layer3_out_311_U.if_empty_n;
    assign fifo_intf_1664.wr_en = AESL_inst_myproject.layer3_out_311_U.if_write & AESL_inst_myproject.layer3_out_311_U.if_full_n;
    assign fifo_intf_1664.fifo_rd_block = 0;
    assign fifo_intf_1664.fifo_wr_block = 0;
    assign fifo_intf_1664.finish = finish;
    csv_file_dump fifo_csv_dumper_1664;
    csv_file_dump cstatus_csv_dumper_1664;
    df_fifo_monitor fifo_monitor_1664;
    df_fifo_intf fifo_intf_1665(clock,reset);
    assign fifo_intf_1665.rd_en = AESL_inst_myproject.layer3_out_312_U.if_read & AESL_inst_myproject.layer3_out_312_U.if_empty_n;
    assign fifo_intf_1665.wr_en = AESL_inst_myproject.layer3_out_312_U.if_write & AESL_inst_myproject.layer3_out_312_U.if_full_n;
    assign fifo_intf_1665.fifo_rd_block = 0;
    assign fifo_intf_1665.fifo_wr_block = 0;
    assign fifo_intf_1665.finish = finish;
    csv_file_dump fifo_csv_dumper_1665;
    csv_file_dump cstatus_csv_dumper_1665;
    df_fifo_monitor fifo_monitor_1665;
    df_fifo_intf fifo_intf_1666(clock,reset);
    assign fifo_intf_1666.rd_en = AESL_inst_myproject.layer3_out_313_U.if_read & AESL_inst_myproject.layer3_out_313_U.if_empty_n;
    assign fifo_intf_1666.wr_en = AESL_inst_myproject.layer3_out_313_U.if_write & AESL_inst_myproject.layer3_out_313_U.if_full_n;
    assign fifo_intf_1666.fifo_rd_block = 0;
    assign fifo_intf_1666.fifo_wr_block = 0;
    assign fifo_intf_1666.finish = finish;
    csv_file_dump fifo_csv_dumper_1666;
    csv_file_dump cstatus_csv_dumper_1666;
    df_fifo_monitor fifo_monitor_1666;
    df_fifo_intf fifo_intf_1667(clock,reset);
    assign fifo_intf_1667.rd_en = AESL_inst_myproject.layer3_out_314_U.if_read & AESL_inst_myproject.layer3_out_314_U.if_empty_n;
    assign fifo_intf_1667.wr_en = AESL_inst_myproject.layer3_out_314_U.if_write & AESL_inst_myproject.layer3_out_314_U.if_full_n;
    assign fifo_intf_1667.fifo_rd_block = 0;
    assign fifo_intf_1667.fifo_wr_block = 0;
    assign fifo_intf_1667.finish = finish;
    csv_file_dump fifo_csv_dumper_1667;
    csv_file_dump cstatus_csv_dumper_1667;
    df_fifo_monitor fifo_monitor_1667;
    df_fifo_intf fifo_intf_1668(clock,reset);
    assign fifo_intf_1668.rd_en = AESL_inst_myproject.layer3_out_315_U.if_read & AESL_inst_myproject.layer3_out_315_U.if_empty_n;
    assign fifo_intf_1668.wr_en = AESL_inst_myproject.layer3_out_315_U.if_write & AESL_inst_myproject.layer3_out_315_U.if_full_n;
    assign fifo_intf_1668.fifo_rd_block = 0;
    assign fifo_intf_1668.fifo_wr_block = 0;
    assign fifo_intf_1668.finish = finish;
    csv_file_dump fifo_csv_dumper_1668;
    csv_file_dump cstatus_csv_dumper_1668;
    df_fifo_monitor fifo_monitor_1668;
    df_fifo_intf fifo_intf_1669(clock,reset);
    assign fifo_intf_1669.rd_en = AESL_inst_myproject.layer3_out_316_U.if_read & AESL_inst_myproject.layer3_out_316_U.if_empty_n;
    assign fifo_intf_1669.wr_en = AESL_inst_myproject.layer3_out_316_U.if_write & AESL_inst_myproject.layer3_out_316_U.if_full_n;
    assign fifo_intf_1669.fifo_rd_block = 0;
    assign fifo_intf_1669.fifo_wr_block = 0;
    assign fifo_intf_1669.finish = finish;
    csv_file_dump fifo_csv_dumper_1669;
    csv_file_dump cstatus_csv_dumper_1669;
    df_fifo_monitor fifo_monitor_1669;
    df_fifo_intf fifo_intf_1670(clock,reset);
    assign fifo_intf_1670.rd_en = AESL_inst_myproject.layer3_out_317_U.if_read & AESL_inst_myproject.layer3_out_317_U.if_empty_n;
    assign fifo_intf_1670.wr_en = AESL_inst_myproject.layer3_out_317_U.if_write & AESL_inst_myproject.layer3_out_317_U.if_full_n;
    assign fifo_intf_1670.fifo_rd_block = 0;
    assign fifo_intf_1670.fifo_wr_block = 0;
    assign fifo_intf_1670.finish = finish;
    csv_file_dump fifo_csv_dumper_1670;
    csv_file_dump cstatus_csv_dumper_1670;
    df_fifo_monitor fifo_monitor_1670;
    df_fifo_intf fifo_intf_1671(clock,reset);
    assign fifo_intf_1671.rd_en = AESL_inst_myproject.layer3_out_318_U.if_read & AESL_inst_myproject.layer3_out_318_U.if_empty_n;
    assign fifo_intf_1671.wr_en = AESL_inst_myproject.layer3_out_318_U.if_write & AESL_inst_myproject.layer3_out_318_U.if_full_n;
    assign fifo_intf_1671.fifo_rd_block = 0;
    assign fifo_intf_1671.fifo_wr_block = 0;
    assign fifo_intf_1671.finish = finish;
    csv_file_dump fifo_csv_dumper_1671;
    csv_file_dump cstatus_csv_dumper_1671;
    df_fifo_monitor fifo_monitor_1671;
    df_fifo_intf fifo_intf_1672(clock,reset);
    assign fifo_intf_1672.rd_en = AESL_inst_myproject.layer3_out_319_U.if_read & AESL_inst_myproject.layer3_out_319_U.if_empty_n;
    assign fifo_intf_1672.wr_en = AESL_inst_myproject.layer3_out_319_U.if_write & AESL_inst_myproject.layer3_out_319_U.if_full_n;
    assign fifo_intf_1672.fifo_rd_block = 0;
    assign fifo_intf_1672.fifo_wr_block = 0;
    assign fifo_intf_1672.finish = finish;
    csv_file_dump fifo_csv_dumper_1672;
    csv_file_dump cstatus_csv_dumper_1672;
    df_fifo_monitor fifo_monitor_1672;
    df_fifo_intf fifo_intf_1673(clock,reset);
    assign fifo_intf_1673.rd_en = AESL_inst_myproject.layer3_out_320_U.if_read & AESL_inst_myproject.layer3_out_320_U.if_empty_n;
    assign fifo_intf_1673.wr_en = AESL_inst_myproject.layer3_out_320_U.if_write & AESL_inst_myproject.layer3_out_320_U.if_full_n;
    assign fifo_intf_1673.fifo_rd_block = 0;
    assign fifo_intf_1673.fifo_wr_block = 0;
    assign fifo_intf_1673.finish = finish;
    csv_file_dump fifo_csv_dumper_1673;
    csv_file_dump cstatus_csv_dumper_1673;
    df_fifo_monitor fifo_monitor_1673;
    df_fifo_intf fifo_intf_1674(clock,reset);
    assign fifo_intf_1674.rd_en = AESL_inst_myproject.layer3_out_321_U.if_read & AESL_inst_myproject.layer3_out_321_U.if_empty_n;
    assign fifo_intf_1674.wr_en = AESL_inst_myproject.layer3_out_321_U.if_write & AESL_inst_myproject.layer3_out_321_U.if_full_n;
    assign fifo_intf_1674.fifo_rd_block = 0;
    assign fifo_intf_1674.fifo_wr_block = 0;
    assign fifo_intf_1674.finish = finish;
    csv_file_dump fifo_csv_dumper_1674;
    csv_file_dump cstatus_csv_dumper_1674;
    df_fifo_monitor fifo_monitor_1674;
    df_fifo_intf fifo_intf_1675(clock,reset);
    assign fifo_intf_1675.rd_en = AESL_inst_myproject.layer3_out_322_U.if_read & AESL_inst_myproject.layer3_out_322_U.if_empty_n;
    assign fifo_intf_1675.wr_en = AESL_inst_myproject.layer3_out_322_U.if_write & AESL_inst_myproject.layer3_out_322_U.if_full_n;
    assign fifo_intf_1675.fifo_rd_block = 0;
    assign fifo_intf_1675.fifo_wr_block = 0;
    assign fifo_intf_1675.finish = finish;
    csv_file_dump fifo_csv_dumper_1675;
    csv_file_dump cstatus_csv_dumper_1675;
    df_fifo_monitor fifo_monitor_1675;
    df_fifo_intf fifo_intf_1676(clock,reset);
    assign fifo_intf_1676.rd_en = AESL_inst_myproject.layer3_out_323_U.if_read & AESL_inst_myproject.layer3_out_323_U.if_empty_n;
    assign fifo_intf_1676.wr_en = AESL_inst_myproject.layer3_out_323_U.if_write & AESL_inst_myproject.layer3_out_323_U.if_full_n;
    assign fifo_intf_1676.fifo_rd_block = 0;
    assign fifo_intf_1676.fifo_wr_block = 0;
    assign fifo_intf_1676.finish = finish;
    csv_file_dump fifo_csv_dumper_1676;
    csv_file_dump cstatus_csv_dumper_1676;
    df_fifo_monitor fifo_monitor_1676;
    df_fifo_intf fifo_intf_1677(clock,reset);
    assign fifo_intf_1677.rd_en = AESL_inst_myproject.layer3_out_324_U.if_read & AESL_inst_myproject.layer3_out_324_U.if_empty_n;
    assign fifo_intf_1677.wr_en = AESL_inst_myproject.layer3_out_324_U.if_write & AESL_inst_myproject.layer3_out_324_U.if_full_n;
    assign fifo_intf_1677.fifo_rd_block = 0;
    assign fifo_intf_1677.fifo_wr_block = 0;
    assign fifo_intf_1677.finish = finish;
    csv_file_dump fifo_csv_dumper_1677;
    csv_file_dump cstatus_csv_dumper_1677;
    df_fifo_monitor fifo_monitor_1677;
    df_fifo_intf fifo_intf_1678(clock,reset);
    assign fifo_intf_1678.rd_en = AESL_inst_myproject.layer3_out_325_U.if_read & AESL_inst_myproject.layer3_out_325_U.if_empty_n;
    assign fifo_intf_1678.wr_en = AESL_inst_myproject.layer3_out_325_U.if_write & AESL_inst_myproject.layer3_out_325_U.if_full_n;
    assign fifo_intf_1678.fifo_rd_block = 0;
    assign fifo_intf_1678.fifo_wr_block = 0;
    assign fifo_intf_1678.finish = finish;
    csv_file_dump fifo_csv_dumper_1678;
    csv_file_dump cstatus_csv_dumper_1678;
    df_fifo_monitor fifo_monitor_1678;
    df_fifo_intf fifo_intf_1679(clock,reset);
    assign fifo_intf_1679.rd_en = AESL_inst_myproject.layer3_out_326_U.if_read & AESL_inst_myproject.layer3_out_326_U.if_empty_n;
    assign fifo_intf_1679.wr_en = AESL_inst_myproject.layer3_out_326_U.if_write & AESL_inst_myproject.layer3_out_326_U.if_full_n;
    assign fifo_intf_1679.fifo_rd_block = 0;
    assign fifo_intf_1679.fifo_wr_block = 0;
    assign fifo_intf_1679.finish = finish;
    csv_file_dump fifo_csv_dumper_1679;
    csv_file_dump cstatus_csv_dumper_1679;
    df_fifo_monitor fifo_monitor_1679;
    df_fifo_intf fifo_intf_1680(clock,reset);
    assign fifo_intf_1680.rd_en = AESL_inst_myproject.layer3_out_327_U.if_read & AESL_inst_myproject.layer3_out_327_U.if_empty_n;
    assign fifo_intf_1680.wr_en = AESL_inst_myproject.layer3_out_327_U.if_write & AESL_inst_myproject.layer3_out_327_U.if_full_n;
    assign fifo_intf_1680.fifo_rd_block = 0;
    assign fifo_intf_1680.fifo_wr_block = 0;
    assign fifo_intf_1680.finish = finish;
    csv_file_dump fifo_csv_dumper_1680;
    csv_file_dump cstatus_csv_dumper_1680;
    df_fifo_monitor fifo_monitor_1680;
    df_fifo_intf fifo_intf_1681(clock,reset);
    assign fifo_intf_1681.rd_en = AESL_inst_myproject.layer3_out_328_U.if_read & AESL_inst_myproject.layer3_out_328_U.if_empty_n;
    assign fifo_intf_1681.wr_en = AESL_inst_myproject.layer3_out_328_U.if_write & AESL_inst_myproject.layer3_out_328_U.if_full_n;
    assign fifo_intf_1681.fifo_rd_block = 0;
    assign fifo_intf_1681.fifo_wr_block = 0;
    assign fifo_intf_1681.finish = finish;
    csv_file_dump fifo_csv_dumper_1681;
    csv_file_dump cstatus_csv_dumper_1681;
    df_fifo_monitor fifo_monitor_1681;
    df_fifo_intf fifo_intf_1682(clock,reset);
    assign fifo_intf_1682.rd_en = AESL_inst_myproject.layer3_out_329_U.if_read & AESL_inst_myproject.layer3_out_329_U.if_empty_n;
    assign fifo_intf_1682.wr_en = AESL_inst_myproject.layer3_out_329_U.if_write & AESL_inst_myproject.layer3_out_329_U.if_full_n;
    assign fifo_intf_1682.fifo_rd_block = 0;
    assign fifo_intf_1682.fifo_wr_block = 0;
    assign fifo_intf_1682.finish = finish;
    csv_file_dump fifo_csv_dumper_1682;
    csv_file_dump cstatus_csv_dumper_1682;
    df_fifo_monitor fifo_monitor_1682;
    df_fifo_intf fifo_intf_1683(clock,reset);
    assign fifo_intf_1683.rd_en = AESL_inst_myproject.layer3_out_330_U.if_read & AESL_inst_myproject.layer3_out_330_U.if_empty_n;
    assign fifo_intf_1683.wr_en = AESL_inst_myproject.layer3_out_330_U.if_write & AESL_inst_myproject.layer3_out_330_U.if_full_n;
    assign fifo_intf_1683.fifo_rd_block = 0;
    assign fifo_intf_1683.fifo_wr_block = 0;
    assign fifo_intf_1683.finish = finish;
    csv_file_dump fifo_csv_dumper_1683;
    csv_file_dump cstatus_csv_dumper_1683;
    df_fifo_monitor fifo_monitor_1683;
    df_fifo_intf fifo_intf_1684(clock,reset);
    assign fifo_intf_1684.rd_en = AESL_inst_myproject.layer3_out_331_U.if_read & AESL_inst_myproject.layer3_out_331_U.if_empty_n;
    assign fifo_intf_1684.wr_en = AESL_inst_myproject.layer3_out_331_U.if_write & AESL_inst_myproject.layer3_out_331_U.if_full_n;
    assign fifo_intf_1684.fifo_rd_block = 0;
    assign fifo_intf_1684.fifo_wr_block = 0;
    assign fifo_intf_1684.finish = finish;
    csv_file_dump fifo_csv_dumper_1684;
    csv_file_dump cstatus_csv_dumper_1684;
    df_fifo_monitor fifo_monitor_1684;
    df_fifo_intf fifo_intf_1685(clock,reset);
    assign fifo_intf_1685.rd_en = AESL_inst_myproject.layer3_out_332_U.if_read & AESL_inst_myproject.layer3_out_332_U.if_empty_n;
    assign fifo_intf_1685.wr_en = AESL_inst_myproject.layer3_out_332_U.if_write & AESL_inst_myproject.layer3_out_332_U.if_full_n;
    assign fifo_intf_1685.fifo_rd_block = 0;
    assign fifo_intf_1685.fifo_wr_block = 0;
    assign fifo_intf_1685.finish = finish;
    csv_file_dump fifo_csv_dumper_1685;
    csv_file_dump cstatus_csv_dumper_1685;
    df_fifo_monitor fifo_monitor_1685;
    df_fifo_intf fifo_intf_1686(clock,reset);
    assign fifo_intf_1686.rd_en = AESL_inst_myproject.layer3_out_333_U.if_read & AESL_inst_myproject.layer3_out_333_U.if_empty_n;
    assign fifo_intf_1686.wr_en = AESL_inst_myproject.layer3_out_333_U.if_write & AESL_inst_myproject.layer3_out_333_U.if_full_n;
    assign fifo_intf_1686.fifo_rd_block = 0;
    assign fifo_intf_1686.fifo_wr_block = 0;
    assign fifo_intf_1686.finish = finish;
    csv_file_dump fifo_csv_dumper_1686;
    csv_file_dump cstatus_csv_dumper_1686;
    df_fifo_monitor fifo_monitor_1686;
    df_fifo_intf fifo_intf_1687(clock,reset);
    assign fifo_intf_1687.rd_en = AESL_inst_myproject.layer3_out_334_U.if_read & AESL_inst_myproject.layer3_out_334_U.if_empty_n;
    assign fifo_intf_1687.wr_en = AESL_inst_myproject.layer3_out_334_U.if_write & AESL_inst_myproject.layer3_out_334_U.if_full_n;
    assign fifo_intf_1687.fifo_rd_block = 0;
    assign fifo_intf_1687.fifo_wr_block = 0;
    assign fifo_intf_1687.finish = finish;
    csv_file_dump fifo_csv_dumper_1687;
    csv_file_dump cstatus_csv_dumper_1687;
    df_fifo_monitor fifo_monitor_1687;
    df_fifo_intf fifo_intf_1688(clock,reset);
    assign fifo_intf_1688.rd_en = AESL_inst_myproject.layer3_out_335_U.if_read & AESL_inst_myproject.layer3_out_335_U.if_empty_n;
    assign fifo_intf_1688.wr_en = AESL_inst_myproject.layer3_out_335_U.if_write & AESL_inst_myproject.layer3_out_335_U.if_full_n;
    assign fifo_intf_1688.fifo_rd_block = 0;
    assign fifo_intf_1688.fifo_wr_block = 0;
    assign fifo_intf_1688.finish = finish;
    csv_file_dump fifo_csv_dumper_1688;
    csv_file_dump cstatus_csv_dumper_1688;
    df_fifo_monitor fifo_monitor_1688;
    df_fifo_intf fifo_intf_1689(clock,reset);
    assign fifo_intf_1689.rd_en = AESL_inst_myproject.layer3_out_336_U.if_read & AESL_inst_myproject.layer3_out_336_U.if_empty_n;
    assign fifo_intf_1689.wr_en = AESL_inst_myproject.layer3_out_336_U.if_write & AESL_inst_myproject.layer3_out_336_U.if_full_n;
    assign fifo_intf_1689.fifo_rd_block = 0;
    assign fifo_intf_1689.fifo_wr_block = 0;
    assign fifo_intf_1689.finish = finish;
    csv_file_dump fifo_csv_dumper_1689;
    csv_file_dump cstatus_csv_dumper_1689;
    df_fifo_monitor fifo_monitor_1689;
    df_fifo_intf fifo_intf_1690(clock,reset);
    assign fifo_intf_1690.rd_en = AESL_inst_myproject.layer3_out_337_U.if_read & AESL_inst_myproject.layer3_out_337_U.if_empty_n;
    assign fifo_intf_1690.wr_en = AESL_inst_myproject.layer3_out_337_U.if_write & AESL_inst_myproject.layer3_out_337_U.if_full_n;
    assign fifo_intf_1690.fifo_rd_block = 0;
    assign fifo_intf_1690.fifo_wr_block = 0;
    assign fifo_intf_1690.finish = finish;
    csv_file_dump fifo_csv_dumper_1690;
    csv_file_dump cstatus_csv_dumper_1690;
    df_fifo_monitor fifo_monitor_1690;
    df_fifo_intf fifo_intf_1691(clock,reset);
    assign fifo_intf_1691.rd_en = AESL_inst_myproject.layer3_out_338_U.if_read & AESL_inst_myproject.layer3_out_338_U.if_empty_n;
    assign fifo_intf_1691.wr_en = AESL_inst_myproject.layer3_out_338_U.if_write & AESL_inst_myproject.layer3_out_338_U.if_full_n;
    assign fifo_intf_1691.fifo_rd_block = 0;
    assign fifo_intf_1691.fifo_wr_block = 0;
    assign fifo_intf_1691.finish = finish;
    csv_file_dump fifo_csv_dumper_1691;
    csv_file_dump cstatus_csv_dumper_1691;
    df_fifo_monitor fifo_monitor_1691;
    df_fifo_intf fifo_intf_1692(clock,reset);
    assign fifo_intf_1692.rd_en = AESL_inst_myproject.layer3_out_339_U.if_read & AESL_inst_myproject.layer3_out_339_U.if_empty_n;
    assign fifo_intf_1692.wr_en = AESL_inst_myproject.layer3_out_339_U.if_write & AESL_inst_myproject.layer3_out_339_U.if_full_n;
    assign fifo_intf_1692.fifo_rd_block = 0;
    assign fifo_intf_1692.fifo_wr_block = 0;
    assign fifo_intf_1692.finish = finish;
    csv_file_dump fifo_csv_dumper_1692;
    csv_file_dump cstatus_csv_dumper_1692;
    df_fifo_monitor fifo_monitor_1692;
    df_fifo_intf fifo_intf_1693(clock,reset);
    assign fifo_intf_1693.rd_en = AESL_inst_myproject.layer3_out_340_U.if_read & AESL_inst_myproject.layer3_out_340_U.if_empty_n;
    assign fifo_intf_1693.wr_en = AESL_inst_myproject.layer3_out_340_U.if_write & AESL_inst_myproject.layer3_out_340_U.if_full_n;
    assign fifo_intf_1693.fifo_rd_block = 0;
    assign fifo_intf_1693.fifo_wr_block = 0;
    assign fifo_intf_1693.finish = finish;
    csv_file_dump fifo_csv_dumper_1693;
    csv_file_dump cstatus_csv_dumper_1693;
    df_fifo_monitor fifo_monitor_1693;
    df_fifo_intf fifo_intf_1694(clock,reset);
    assign fifo_intf_1694.rd_en = AESL_inst_myproject.layer3_out_341_U.if_read & AESL_inst_myproject.layer3_out_341_U.if_empty_n;
    assign fifo_intf_1694.wr_en = AESL_inst_myproject.layer3_out_341_U.if_write & AESL_inst_myproject.layer3_out_341_U.if_full_n;
    assign fifo_intf_1694.fifo_rd_block = 0;
    assign fifo_intf_1694.fifo_wr_block = 0;
    assign fifo_intf_1694.finish = finish;
    csv_file_dump fifo_csv_dumper_1694;
    csv_file_dump cstatus_csv_dumper_1694;
    df_fifo_monitor fifo_monitor_1694;
    df_fifo_intf fifo_intf_1695(clock,reset);
    assign fifo_intf_1695.rd_en = AESL_inst_myproject.layer3_out_342_U.if_read & AESL_inst_myproject.layer3_out_342_U.if_empty_n;
    assign fifo_intf_1695.wr_en = AESL_inst_myproject.layer3_out_342_U.if_write & AESL_inst_myproject.layer3_out_342_U.if_full_n;
    assign fifo_intf_1695.fifo_rd_block = 0;
    assign fifo_intf_1695.fifo_wr_block = 0;
    assign fifo_intf_1695.finish = finish;
    csv_file_dump fifo_csv_dumper_1695;
    csv_file_dump cstatus_csv_dumper_1695;
    df_fifo_monitor fifo_monitor_1695;
    df_fifo_intf fifo_intf_1696(clock,reset);
    assign fifo_intf_1696.rd_en = AESL_inst_myproject.layer3_out_343_U.if_read & AESL_inst_myproject.layer3_out_343_U.if_empty_n;
    assign fifo_intf_1696.wr_en = AESL_inst_myproject.layer3_out_343_U.if_write & AESL_inst_myproject.layer3_out_343_U.if_full_n;
    assign fifo_intf_1696.fifo_rd_block = 0;
    assign fifo_intf_1696.fifo_wr_block = 0;
    assign fifo_intf_1696.finish = finish;
    csv_file_dump fifo_csv_dumper_1696;
    csv_file_dump cstatus_csv_dumper_1696;
    df_fifo_monitor fifo_monitor_1696;
    df_fifo_intf fifo_intf_1697(clock,reset);
    assign fifo_intf_1697.rd_en = AESL_inst_myproject.layer3_out_344_U.if_read & AESL_inst_myproject.layer3_out_344_U.if_empty_n;
    assign fifo_intf_1697.wr_en = AESL_inst_myproject.layer3_out_344_U.if_write & AESL_inst_myproject.layer3_out_344_U.if_full_n;
    assign fifo_intf_1697.fifo_rd_block = 0;
    assign fifo_intf_1697.fifo_wr_block = 0;
    assign fifo_intf_1697.finish = finish;
    csv_file_dump fifo_csv_dumper_1697;
    csv_file_dump cstatus_csv_dumper_1697;
    df_fifo_monitor fifo_monitor_1697;
    df_fifo_intf fifo_intf_1698(clock,reset);
    assign fifo_intf_1698.rd_en = AESL_inst_myproject.layer3_out_345_U.if_read & AESL_inst_myproject.layer3_out_345_U.if_empty_n;
    assign fifo_intf_1698.wr_en = AESL_inst_myproject.layer3_out_345_U.if_write & AESL_inst_myproject.layer3_out_345_U.if_full_n;
    assign fifo_intf_1698.fifo_rd_block = 0;
    assign fifo_intf_1698.fifo_wr_block = 0;
    assign fifo_intf_1698.finish = finish;
    csv_file_dump fifo_csv_dumper_1698;
    csv_file_dump cstatus_csv_dumper_1698;
    df_fifo_monitor fifo_monitor_1698;
    df_fifo_intf fifo_intf_1699(clock,reset);
    assign fifo_intf_1699.rd_en = AESL_inst_myproject.layer3_out_346_U.if_read & AESL_inst_myproject.layer3_out_346_U.if_empty_n;
    assign fifo_intf_1699.wr_en = AESL_inst_myproject.layer3_out_346_U.if_write & AESL_inst_myproject.layer3_out_346_U.if_full_n;
    assign fifo_intf_1699.fifo_rd_block = 0;
    assign fifo_intf_1699.fifo_wr_block = 0;
    assign fifo_intf_1699.finish = finish;
    csv_file_dump fifo_csv_dumper_1699;
    csv_file_dump cstatus_csv_dumper_1699;
    df_fifo_monitor fifo_monitor_1699;
    df_fifo_intf fifo_intf_1700(clock,reset);
    assign fifo_intf_1700.rd_en = AESL_inst_myproject.layer3_out_347_U.if_read & AESL_inst_myproject.layer3_out_347_U.if_empty_n;
    assign fifo_intf_1700.wr_en = AESL_inst_myproject.layer3_out_347_U.if_write & AESL_inst_myproject.layer3_out_347_U.if_full_n;
    assign fifo_intf_1700.fifo_rd_block = 0;
    assign fifo_intf_1700.fifo_wr_block = 0;
    assign fifo_intf_1700.finish = finish;
    csv_file_dump fifo_csv_dumper_1700;
    csv_file_dump cstatus_csv_dumper_1700;
    df_fifo_monitor fifo_monitor_1700;
    df_fifo_intf fifo_intf_1701(clock,reset);
    assign fifo_intf_1701.rd_en = AESL_inst_myproject.layer3_out_348_U.if_read & AESL_inst_myproject.layer3_out_348_U.if_empty_n;
    assign fifo_intf_1701.wr_en = AESL_inst_myproject.layer3_out_348_U.if_write & AESL_inst_myproject.layer3_out_348_U.if_full_n;
    assign fifo_intf_1701.fifo_rd_block = 0;
    assign fifo_intf_1701.fifo_wr_block = 0;
    assign fifo_intf_1701.finish = finish;
    csv_file_dump fifo_csv_dumper_1701;
    csv_file_dump cstatus_csv_dumper_1701;
    df_fifo_monitor fifo_monitor_1701;
    df_fifo_intf fifo_intf_1702(clock,reset);
    assign fifo_intf_1702.rd_en = AESL_inst_myproject.layer3_out_349_U.if_read & AESL_inst_myproject.layer3_out_349_U.if_empty_n;
    assign fifo_intf_1702.wr_en = AESL_inst_myproject.layer3_out_349_U.if_write & AESL_inst_myproject.layer3_out_349_U.if_full_n;
    assign fifo_intf_1702.fifo_rd_block = 0;
    assign fifo_intf_1702.fifo_wr_block = 0;
    assign fifo_intf_1702.finish = finish;
    csv_file_dump fifo_csv_dumper_1702;
    csv_file_dump cstatus_csv_dumper_1702;
    df_fifo_monitor fifo_monitor_1702;
    df_fifo_intf fifo_intf_1703(clock,reset);
    assign fifo_intf_1703.rd_en = AESL_inst_myproject.layer3_out_350_U.if_read & AESL_inst_myproject.layer3_out_350_U.if_empty_n;
    assign fifo_intf_1703.wr_en = AESL_inst_myproject.layer3_out_350_U.if_write & AESL_inst_myproject.layer3_out_350_U.if_full_n;
    assign fifo_intf_1703.fifo_rd_block = 0;
    assign fifo_intf_1703.fifo_wr_block = 0;
    assign fifo_intf_1703.finish = finish;
    csv_file_dump fifo_csv_dumper_1703;
    csv_file_dump cstatus_csv_dumper_1703;
    df_fifo_monitor fifo_monitor_1703;
    df_fifo_intf fifo_intf_1704(clock,reset);
    assign fifo_intf_1704.rd_en = AESL_inst_myproject.layer3_out_351_U.if_read & AESL_inst_myproject.layer3_out_351_U.if_empty_n;
    assign fifo_intf_1704.wr_en = AESL_inst_myproject.layer3_out_351_U.if_write & AESL_inst_myproject.layer3_out_351_U.if_full_n;
    assign fifo_intf_1704.fifo_rd_block = 0;
    assign fifo_intf_1704.fifo_wr_block = 0;
    assign fifo_intf_1704.finish = finish;
    csv_file_dump fifo_csv_dumper_1704;
    csv_file_dump cstatus_csv_dumper_1704;
    df_fifo_monitor fifo_monitor_1704;
    df_fifo_intf fifo_intf_1705(clock,reset);
    assign fifo_intf_1705.rd_en = AESL_inst_myproject.layer3_out_352_U.if_read & AESL_inst_myproject.layer3_out_352_U.if_empty_n;
    assign fifo_intf_1705.wr_en = AESL_inst_myproject.layer3_out_352_U.if_write & AESL_inst_myproject.layer3_out_352_U.if_full_n;
    assign fifo_intf_1705.fifo_rd_block = 0;
    assign fifo_intf_1705.fifo_wr_block = 0;
    assign fifo_intf_1705.finish = finish;
    csv_file_dump fifo_csv_dumper_1705;
    csv_file_dump cstatus_csv_dumper_1705;
    df_fifo_monitor fifo_monitor_1705;
    df_fifo_intf fifo_intf_1706(clock,reset);
    assign fifo_intf_1706.rd_en = AESL_inst_myproject.layer3_out_353_U.if_read & AESL_inst_myproject.layer3_out_353_U.if_empty_n;
    assign fifo_intf_1706.wr_en = AESL_inst_myproject.layer3_out_353_U.if_write & AESL_inst_myproject.layer3_out_353_U.if_full_n;
    assign fifo_intf_1706.fifo_rd_block = 0;
    assign fifo_intf_1706.fifo_wr_block = 0;
    assign fifo_intf_1706.finish = finish;
    csv_file_dump fifo_csv_dumper_1706;
    csv_file_dump cstatus_csv_dumper_1706;
    df_fifo_monitor fifo_monitor_1706;
    df_fifo_intf fifo_intf_1707(clock,reset);
    assign fifo_intf_1707.rd_en = AESL_inst_myproject.layer3_out_354_U.if_read & AESL_inst_myproject.layer3_out_354_U.if_empty_n;
    assign fifo_intf_1707.wr_en = AESL_inst_myproject.layer3_out_354_U.if_write & AESL_inst_myproject.layer3_out_354_U.if_full_n;
    assign fifo_intf_1707.fifo_rd_block = 0;
    assign fifo_intf_1707.fifo_wr_block = 0;
    assign fifo_intf_1707.finish = finish;
    csv_file_dump fifo_csv_dumper_1707;
    csv_file_dump cstatus_csv_dumper_1707;
    df_fifo_monitor fifo_monitor_1707;
    df_fifo_intf fifo_intf_1708(clock,reset);
    assign fifo_intf_1708.rd_en = AESL_inst_myproject.layer3_out_355_U.if_read & AESL_inst_myproject.layer3_out_355_U.if_empty_n;
    assign fifo_intf_1708.wr_en = AESL_inst_myproject.layer3_out_355_U.if_write & AESL_inst_myproject.layer3_out_355_U.if_full_n;
    assign fifo_intf_1708.fifo_rd_block = 0;
    assign fifo_intf_1708.fifo_wr_block = 0;
    assign fifo_intf_1708.finish = finish;
    csv_file_dump fifo_csv_dumper_1708;
    csv_file_dump cstatus_csv_dumper_1708;
    df_fifo_monitor fifo_monitor_1708;
    df_fifo_intf fifo_intf_1709(clock,reset);
    assign fifo_intf_1709.rd_en = AESL_inst_myproject.layer3_out_356_U.if_read & AESL_inst_myproject.layer3_out_356_U.if_empty_n;
    assign fifo_intf_1709.wr_en = AESL_inst_myproject.layer3_out_356_U.if_write & AESL_inst_myproject.layer3_out_356_U.if_full_n;
    assign fifo_intf_1709.fifo_rd_block = 0;
    assign fifo_intf_1709.fifo_wr_block = 0;
    assign fifo_intf_1709.finish = finish;
    csv_file_dump fifo_csv_dumper_1709;
    csv_file_dump cstatus_csv_dumper_1709;
    df_fifo_monitor fifo_monitor_1709;
    df_fifo_intf fifo_intf_1710(clock,reset);
    assign fifo_intf_1710.rd_en = AESL_inst_myproject.layer3_out_357_U.if_read & AESL_inst_myproject.layer3_out_357_U.if_empty_n;
    assign fifo_intf_1710.wr_en = AESL_inst_myproject.layer3_out_357_U.if_write & AESL_inst_myproject.layer3_out_357_U.if_full_n;
    assign fifo_intf_1710.fifo_rd_block = 0;
    assign fifo_intf_1710.fifo_wr_block = 0;
    assign fifo_intf_1710.finish = finish;
    csv_file_dump fifo_csv_dumper_1710;
    csv_file_dump cstatus_csv_dumper_1710;
    df_fifo_monitor fifo_monitor_1710;
    df_fifo_intf fifo_intf_1711(clock,reset);
    assign fifo_intf_1711.rd_en = AESL_inst_myproject.layer3_out_358_U.if_read & AESL_inst_myproject.layer3_out_358_U.if_empty_n;
    assign fifo_intf_1711.wr_en = AESL_inst_myproject.layer3_out_358_U.if_write & AESL_inst_myproject.layer3_out_358_U.if_full_n;
    assign fifo_intf_1711.fifo_rd_block = 0;
    assign fifo_intf_1711.fifo_wr_block = 0;
    assign fifo_intf_1711.finish = finish;
    csv_file_dump fifo_csv_dumper_1711;
    csv_file_dump cstatus_csv_dumper_1711;
    df_fifo_monitor fifo_monitor_1711;
    df_fifo_intf fifo_intf_1712(clock,reset);
    assign fifo_intf_1712.rd_en = AESL_inst_myproject.layer3_out_359_U.if_read & AESL_inst_myproject.layer3_out_359_U.if_empty_n;
    assign fifo_intf_1712.wr_en = AESL_inst_myproject.layer3_out_359_U.if_write & AESL_inst_myproject.layer3_out_359_U.if_full_n;
    assign fifo_intf_1712.fifo_rd_block = 0;
    assign fifo_intf_1712.fifo_wr_block = 0;
    assign fifo_intf_1712.finish = finish;
    csv_file_dump fifo_csv_dumper_1712;
    csv_file_dump cstatus_csv_dumper_1712;
    df_fifo_monitor fifo_monitor_1712;
    df_fifo_intf fifo_intf_1713(clock,reset);
    assign fifo_intf_1713.rd_en = AESL_inst_myproject.layer3_out_360_U.if_read & AESL_inst_myproject.layer3_out_360_U.if_empty_n;
    assign fifo_intf_1713.wr_en = AESL_inst_myproject.layer3_out_360_U.if_write & AESL_inst_myproject.layer3_out_360_U.if_full_n;
    assign fifo_intf_1713.fifo_rd_block = 0;
    assign fifo_intf_1713.fifo_wr_block = 0;
    assign fifo_intf_1713.finish = finish;
    csv_file_dump fifo_csv_dumper_1713;
    csv_file_dump cstatus_csv_dumper_1713;
    df_fifo_monitor fifo_monitor_1713;
    df_fifo_intf fifo_intf_1714(clock,reset);
    assign fifo_intf_1714.rd_en = AESL_inst_myproject.layer3_out_361_U.if_read & AESL_inst_myproject.layer3_out_361_U.if_empty_n;
    assign fifo_intf_1714.wr_en = AESL_inst_myproject.layer3_out_361_U.if_write & AESL_inst_myproject.layer3_out_361_U.if_full_n;
    assign fifo_intf_1714.fifo_rd_block = 0;
    assign fifo_intf_1714.fifo_wr_block = 0;
    assign fifo_intf_1714.finish = finish;
    csv_file_dump fifo_csv_dumper_1714;
    csv_file_dump cstatus_csv_dumper_1714;
    df_fifo_monitor fifo_monitor_1714;
    df_fifo_intf fifo_intf_1715(clock,reset);
    assign fifo_intf_1715.rd_en = AESL_inst_myproject.layer3_out_362_U.if_read & AESL_inst_myproject.layer3_out_362_U.if_empty_n;
    assign fifo_intf_1715.wr_en = AESL_inst_myproject.layer3_out_362_U.if_write & AESL_inst_myproject.layer3_out_362_U.if_full_n;
    assign fifo_intf_1715.fifo_rd_block = 0;
    assign fifo_intf_1715.fifo_wr_block = 0;
    assign fifo_intf_1715.finish = finish;
    csv_file_dump fifo_csv_dumper_1715;
    csv_file_dump cstatus_csv_dumper_1715;
    df_fifo_monitor fifo_monitor_1715;
    df_fifo_intf fifo_intf_1716(clock,reset);
    assign fifo_intf_1716.rd_en = AESL_inst_myproject.layer3_out_363_U.if_read & AESL_inst_myproject.layer3_out_363_U.if_empty_n;
    assign fifo_intf_1716.wr_en = AESL_inst_myproject.layer3_out_363_U.if_write & AESL_inst_myproject.layer3_out_363_U.if_full_n;
    assign fifo_intf_1716.fifo_rd_block = 0;
    assign fifo_intf_1716.fifo_wr_block = 0;
    assign fifo_intf_1716.finish = finish;
    csv_file_dump fifo_csv_dumper_1716;
    csv_file_dump cstatus_csv_dumper_1716;
    df_fifo_monitor fifo_monitor_1716;
    df_fifo_intf fifo_intf_1717(clock,reset);
    assign fifo_intf_1717.rd_en = AESL_inst_myproject.layer3_out_364_U.if_read & AESL_inst_myproject.layer3_out_364_U.if_empty_n;
    assign fifo_intf_1717.wr_en = AESL_inst_myproject.layer3_out_364_U.if_write & AESL_inst_myproject.layer3_out_364_U.if_full_n;
    assign fifo_intf_1717.fifo_rd_block = 0;
    assign fifo_intf_1717.fifo_wr_block = 0;
    assign fifo_intf_1717.finish = finish;
    csv_file_dump fifo_csv_dumper_1717;
    csv_file_dump cstatus_csv_dumper_1717;
    df_fifo_monitor fifo_monitor_1717;
    df_fifo_intf fifo_intf_1718(clock,reset);
    assign fifo_intf_1718.rd_en = AESL_inst_myproject.layer3_out_365_U.if_read & AESL_inst_myproject.layer3_out_365_U.if_empty_n;
    assign fifo_intf_1718.wr_en = AESL_inst_myproject.layer3_out_365_U.if_write & AESL_inst_myproject.layer3_out_365_U.if_full_n;
    assign fifo_intf_1718.fifo_rd_block = 0;
    assign fifo_intf_1718.fifo_wr_block = 0;
    assign fifo_intf_1718.finish = finish;
    csv_file_dump fifo_csv_dumper_1718;
    csv_file_dump cstatus_csv_dumper_1718;
    df_fifo_monitor fifo_monitor_1718;
    df_fifo_intf fifo_intf_1719(clock,reset);
    assign fifo_intf_1719.rd_en = AESL_inst_myproject.layer3_out_366_U.if_read & AESL_inst_myproject.layer3_out_366_U.if_empty_n;
    assign fifo_intf_1719.wr_en = AESL_inst_myproject.layer3_out_366_U.if_write & AESL_inst_myproject.layer3_out_366_U.if_full_n;
    assign fifo_intf_1719.fifo_rd_block = 0;
    assign fifo_intf_1719.fifo_wr_block = 0;
    assign fifo_intf_1719.finish = finish;
    csv_file_dump fifo_csv_dumper_1719;
    csv_file_dump cstatus_csv_dumper_1719;
    df_fifo_monitor fifo_monitor_1719;
    df_fifo_intf fifo_intf_1720(clock,reset);
    assign fifo_intf_1720.rd_en = AESL_inst_myproject.layer3_out_367_U.if_read & AESL_inst_myproject.layer3_out_367_U.if_empty_n;
    assign fifo_intf_1720.wr_en = AESL_inst_myproject.layer3_out_367_U.if_write & AESL_inst_myproject.layer3_out_367_U.if_full_n;
    assign fifo_intf_1720.fifo_rd_block = 0;
    assign fifo_intf_1720.fifo_wr_block = 0;
    assign fifo_intf_1720.finish = finish;
    csv_file_dump fifo_csv_dumper_1720;
    csv_file_dump cstatus_csv_dumper_1720;
    df_fifo_monitor fifo_monitor_1720;
    df_fifo_intf fifo_intf_1721(clock,reset);
    assign fifo_intf_1721.rd_en = AESL_inst_myproject.layer3_out_368_U.if_read & AESL_inst_myproject.layer3_out_368_U.if_empty_n;
    assign fifo_intf_1721.wr_en = AESL_inst_myproject.layer3_out_368_U.if_write & AESL_inst_myproject.layer3_out_368_U.if_full_n;
    assign fifo_intf_1721.fifo_rd_block = 0;
    assign fifo_intf_1721.fifo_wr_block = 0;
    assign fifo_intf_1721.finish = finish;
    csv_file_dump fifo_csv_dumper_1721;
    csv_file_dump cstatus_csv_dumper_1721;
    df_fifo_monitor fifo_monitor_1721;
    df_fifo_intf fifo_intf_1722(clock,reset);
    assign fifo_intf_1722.rd_en = AESL_inst_myproject.layer3_out_369_U.if_read & AESL_inst_myproject.layer3_out_369_U.if_empty_n;
    assign fifo_intf_1722.wr_en = AESL_inst_myproject.layer3_out_369_U.if_write & AESL_inst_myproject.layer3_out_369_U.if_full_n;
    assign fifo_intf_1722.fifo_rd_block = 0;
    assign fifo_intf_1722.fifo_wr_block = 0;
    assign fifo_intf_1722.finish = finish;
    csv_file_dump fifo_csv_dumper_1722;
    csv_file_dump cstatus_csv_dumper_1722;
    df_fifo_monitor fifo_monitor_1722;
    df_fifo_intf fifo_intf_1723(clock,reset);
    assign fifo_intf_1723.rd_en = AESL_inst_myproject.layer3_out_370_U.if_read & AESL_inst_myproject.layer3_out_370_U.if_empty_n;
    assign fifo_intf_1723.wr_en = AESL_inst_myproject.layer3_out_370_U.if_write & AESL_inst_myproject.layer3_out_370_U.if_full_n;
    assign fifo_intf_1723.fifo_rd_block = 0;
    assign fifo_intf_1723.fifo_wr_block = 0;
    assign fifo_intf_1723.finish = finish;
    csv_file_dump fifo_csv_dumper_1723;
    csv_file_dump cstatus_csv_dumper_1723;
    df_fifo_monitor fifo_monitor_1723;
    df_fifo_intf fifo_intf_1724(clock,reset);
    assign fifo_intf_1724.rd_en = AESL_inst_myproject.layer3_out_371_U.if_read & AESL_inst_myproject.layer3_out_371_U.if_empty_n;
    assign fifo_intf_1724.wr_en = AESL_inst_myproject.layer3_out_371_U.if_write & AESL_inst_myproject.layer3_out_371_U.if_full_n;
    assign fifo_intf_1724.fifo_rd_block = 0;
    assign fifo_intf_1724.fifo_wr_block = 0;
    assign fifo_intf_1724.finish = finish;
    csv_file_dump fifo_csv_dumper_1724;
    csv_file_dump cstatus_csv_dumper_1724;
    df_fifo_monitor fifo_monitor_1724;
    df_fifo_intf fifo_intf_1725(clock,reset);
    assign fifo_intf_1725.rd_en = AESL_inst_myproject.layer3_out_372_U.if_read & AESL_inst_myproject.layer3_out_372_U.if_empty_n;
    assign fifo_intf_1725.wr_en = AESL_inst_myproject.layer3_out_372_U.if_write & AESL_inst_myproject.layer3_out_372_U.if_full_n;
    assign fifo_intf_1725.fifo_rd_block = 0;
    assign fifo_intf_1725.fifo_wr_block = 0;
    assign fifo_intf_1725.finish = finish;
    csv_file_dump fifo_csv_dumper_1725;
    csv_file_dump cstatus_csv_dumper_1725;
    df_fifo_monitor fifo_monitor_1725;
    df_fifo_intf fifo_intf_1726(clock,reset);
    assign fifo_intf_1726.rd_en = AESL_inst_myproject.layer3_out_373_U.if_read & AESL_inst_myproject.layer3_out_373_U.if_empty_n;
    assign fifo_intf_1726.wr_en = AESL_inst_myproject.layer3_out_373_U.if_write & AESL_inst_myproject.layer3_out_373_U.if_full_n;
    assign fifo_intf_1726.fifo_rd_block = 0;
    assign fifo_intf_1726.fifo_wr_block = 0;
    assign fifo_intf_1726.finish = finish;
    csv_file_dump fifo_csv_dumper_1726;
    csv_file_dump cstatus_csv_dumper_1726;
    df_fifo_monitor fifo_monitor_1726;
    df_fifo_intf fifo_intf_1727(clock,reset);
    assign fifo_intf_1727.rd_en = AESL_inst_myproject.layer3_out_374_U.if_read & AESL_inst_myproject.layer3_out_374_U.if_empty_n;
    assign fifo_intf_1727.wr_en = AESL_inst_myproject.layer3_out_374_U.if_write & AESL_inst_myproject.layer3_out_374_U.if_full_n;
    assign fifo_intf_1727.fifo_rd_block = 0;
    assign fifo_intf_1727.fifo_wr_block = 0;
    assign fifo_intf_1727.finish = finish;
    csv_file_dump fifo_csv_dumper_1727;
    csv_file_dump cstatus_csv_dumper_1727;
    df_fifo_monitor fifo_monitor_1727;
    df_fifo_intf fifo_intf_1728(clock,reset);
    assign fifo_intf_1728.rd_en = AESL_inst_myproject.layer3_out_375_U.if_read & AESL_inst_myproject.layer3_out_375_U.if_empty_n;
    assign fifo_intf_1728.wr_en = AESL_inst_myproject.layer3_out_375_U.if_write & AESL_inst_myproject.layer3_out_375_U.if_full_n;
    assign fifo_intf_1728.fifo_rd_block = 0;
    assign fifo_intf_1728.fifo_wr_block = 0;
    assign fifo_intf_1728.finish = finish;
    csv_file_dump fifo_csv_dumper_1728;
    csv_file_dump cstatus_csv_dumper_1728;
    df_fifo_monitor fifo_monitor_1728;
    df_fifo_intf fifo_intf_1729(clock,reset);
    assign fifo_intf_1729.rd_en = AESL_inst_myproject.layer3_out_376_U.if_read & AESL_inst_myproject.layer3_out_376_U.if_empty_n;
    assign fifo_intf_1729.wr_en = AESL_inst_myproject.layer3_out_376_U.if_write & AESL_inst_myproject.layer3_out_376_U.if_full_n;
    assign fifo_intf_1729.fifo_rd_block = 0;
    assign fifo_intf_1729.fifo_wr_block = 0;
    assign fifo_intf_1729.finish = finish;
    csv_file_dump fifo_csv_dumper_1729;
    csv_file_dump cstatus_csv_dumper_1729;
    df_fifo_monitor fifo_monitor_1729;
    df_fifo_intf fifo_intf_1730(clock,reset);
    assign fifo_intf_1730.rd_en = AESL_inst_myproject.layer3_out_377_U.if_read & AESL_inst_myproject.layer3_out_377_U.if_empty_n;
    assign fifo_intf_1730.wr_en = AESL_inst_myproject.layer3_out_377_U.if_write & AESL_inst_myproject.layer3_out_377_U.if_full_n;
    assign fifo_intf_1730.fifo_rd_block = 0;
    assign fifo_intf_1730.fifo_wr_block = 0;
    assign fifo_intf_1730.finish = finish;
    csv_file_dump fifo_csv_dumper_1730;
    csv_file_dump cstatus_csv_dumper_1730;
    df_fifo_monitor fifo_monitor_1730;
    df_fifo_intf fifo_intf_1731(clock,reset);
    assign fifo_intf_1731.rd_en = AESL_inst_myproject.layer3_out_378_U.if_read & AESL_inst_myproject.layer3_out_378_U.if_empty_n;
    assign fifo_intf_1731.wr_en = AESL_inst_myproject.layer3_out_378_U.if_write & AESL_inst_myproject.layer3_out_378_U.if_full_n;
    assign fifo_intf_1731.fifo_rd_block = 0;
    assign fifo_intf_1731.fifo_wr_block = 0;
    assign fifo_intf_1731.finish = finish;
    csv_file_dump fifo_csv_dumper_1731;
    csv_file_dump cstatus_csv_dumper_1731;
    df_fifo_monitor fifo_monitor_1731;
    df_fifo_intf fifo_intf_1732(clock,reset);
    assign fifo_intf_1732.rd_en = AESL_inst_myproject.layer3_out_379_U.if_read & AESL_inst_myproject.layer3_out_379_U.if_empty_n;
    assign fifo_intf_1732.wr_en = AESL_inst_myproject.layer3_out_379_U.if_write & AESL_inst_myproject.layer3_out_379_U.if_full_n;
    assign fifo_intf_1732.fifo_rd_block = 0;
    assign fifo_intf_1732.fifo_wr_block = 0;
    assign fifo_intf_1732.finish = finish;
    csv_file_dump fifo_csv_dumper_1732;
    csv_file_dump cstatus_csv_dumper_1732;
    df_fifo_monitor fifo_monitor_1732;
    df_fifo_intf fifo_intf_1733(clock,reset);
    assign fifo_intf_1733.rd_en = AESL_inst_myproject.layer3_out_380_U.if_read & AESL_inst_myproject.layer3_out_380_U.if_empty_n;
    assign fifo_intf_1733.wr_en = AESL_inst_myproject.layer3_out_380_U.if_write & AESL_inst_myproject.layer3_out_380_U.if_full_n;
    assign fifo_intf_1733.fifo_rd_block = 0;
    assign fifo_intf_1733.fifo_wr_block = 0;
    assign fifo_intf_1733.finish = finish;
    csv_file_dump fifo_csv_dumper_1733;
    csv_file_dump cstatus_csv_dumper_1733;
    df_fifo_monitor fifo_monitor_1733;
    df_fifo_intf fifo_intf_1734(clock,reset);
    assign fifo_intf_1734.rd_en = AESL_inst_myproject.layer3_out_381_U.if_read & AESL_inst_myproject.layer3_out_381_U.if_empty_n;
    assign fifo_intf_1734.wr_en = AESL_inst_myproject.layer3_out_381_U.if_write & AESL_inst_myproject.layer3_out_381_U.if_full_n;
    assign fifo_intf_1734.fifo_rd_block = 0;
    assign fifo_intf_1734.fifo_wr_block = 0;
    assign fifo_intf_1734.finish = finish;
    csv_file_dump fifo_csv_dumper_1734;
    csv_file_dump cstatus_csv_dumper_1734;
    df_fifo_monitor fifo_monitor_1734;
    df_fifo_intf fifo_intf_1735(clock,reset);
    assign fifo_intf_1735.rd_en = AESL_inst_myproject.layer3_out_382_U.if_read & AESL_inst_myproject.layer3_out_382_U.if_empty_n;
    assign fifo_intf_1735.wr_en = AESL_inst_myproject.layer3_out_382_U.if_write & AESL_inst_myproject.layer3_out_382_U.if_full_n;
    assign fifo_intf_1735.fifo_rd_block = 0;
    assign fifo_intf_1735.fifo_wr_block = 0;
    assign fifo_intf_1735.finish = finish;
    csv_file_dump fifo_csv_dumper_1735;
    csv_file_dump cstatus_csv_dumper_1735;
    df_fifo_monitor fifo_monitor_1735;
    df_fifo_intf fifo_intf_1736(clock,reset);
    assign fifo_intf_1736.rd_en = AESL_inst_myproject.layer3_out_383_U.if_read & AESL_inst_myproject.layer3_out_383_U.if_empty_n;
    assign fifo_intf_1736.wr_en = AESL_inst_myproject.layer3_out_383_U.if_write & AESL_inst_myproject.layer3_out_383_U.if_full_n;
    assign fifo_intf_1736.fifo_rd_block = 0;
    assign fifo_intf_1736.fifo_wr_block = 0;
    assign fifo_intf_1736.finish = finish;
    csv_file_dump fifo_csv_dumper_1736;
    csv_file_dump cstatus_csv_dumper_1736;
    df_fifo_monitor fifo_monitor_1736;
    df_fifo_intf fifo_intf_1737(clock,reset);
    assign fifo_intf_1737.rd_en = AESL_inst_myproject.layer3_out_384_U.if_read & AESL_inst_myproject.layer3_out_384_U.if_empty_n;
    assign fifo_intf_1737.wr_en = AESL_inst_myproject.layer3_out_384_U.if_write & AESL_inst_myproject.layer3_out_384_U.if_full_n;
    assign fifo_intf_1737.fifo_rd_block = 0;
    assign fifo_intf_1737.fifo_wr_block = 0;
    assign fifo_intf_1737.finish = finish;
    csv_file_dump fifo_csv_dumper_1737;
    csv_file_dump cstatus_csv_dumper_1737;
    df_fifo_monitor fifo_monitor_1737;
    df_fifo_intf fifo_intf_1738(clock,reset);
    assign fifo_intf_1738.rd_en = AESL_inst_myproject.layer3_out_385_U.if_read & AESL_inst_myproject.layer3_out_385_U.if_empty_n;
    assign fifo_intf_1738.wr_en = AESL_inst_myproject.layer3_out_385_U.if_write & AESL_inst_myproject.layer3_out_385_U.if_full_n;
    assign fifo_intf_1738.fifo_rd_block = 0;
    assign fifo_intf_1738.fifo_wr_block = 0;
    assign fifo_intf_1738.finish = finish;
    csv_file_dump fifo_csv_dumper_1738;
    csv_file_dump cstatus_csv_dumper_1738;
    df_fifo_monitor fifo_monitor_1738;
    df_fifo_intf fifo_intf_1739(clock,reset);
    assign fifo_intf_1739.rd_en = AESL_inst_myproject.layer3_out_386_U.if_read & AESL_inst_myproject.layer3_out_386_U.if_empty_n;
    assign fifo_intf_1739.wr_en = AESL_inst_myproject.layer3_out_386_U.if_write & AESL_inst_myproject.layer3_out_386_U.if_full_n;
    assign fifo_intf_1739.fifo_rd_block = 0;
    assign fifo_intf_1739.fifo_wr_block = 0;
    assign fifo_intf_1739.finish = finish;
    csv_file_dump fifo_csv_dumper_1739;
    csv_file_dump cstatus_csv_dumper_1739;
    df_fifo_monitor fifo_monitor_1739;
    df_fifo_intf fifo_intf_1740(clock,reset);
    assign fifo_intf_1740.rd_en = AESL_inst_myproject.layer3_out_387_U.if_read & AESL_inst_myproject.layer3_out_387_U.if_empty_n;
    assign fifo_intf_1740.wr_en = AESL_inst_myproject.layer3_out_387_U.if_write & AESL_inst_myproject.layer3_out_387_U.if_full_n;
    assign fifo_intf_1740.fifo_rd_block = 0;
    assign fifo_intf_1740.fifo_wr_block = 0;
    assign fifo_intf_1740.finish = finish;
    csv_file_dump fifo_csv_dumper_1740;
    csv_file_dump cstatus_csv_dumper_1740;
    df_fifo_monitor fifo_monitor_1740;
    df_fifo_intf fifo_intf_1741(clock,reset);
    assign fifo_intf_1741.rd_en = AESL_inst_myproject.layer3_out_388_U.if_read & AESL_inst_myproject.layer3_out_388_U.if_empty_n;
    assign fifo_intf_1741.wr_en = AESL_inst_myproject.layer3_out_388_U.if_write & AESL_inst_myproject.layer3_out_388_U.if_full_n;
    assign fifo_intf_1741.fifo_rd_block = 0;
    assign fifo_intf_1741.fifo_wr_block = 0;
    assign fifo_intf_1741.finish = finish;
    csv_file_dump fifo_csv_dumper_1741;
    csv_file_dump cstatus_csv_dumper_1741;
    df_fifo_monitor fifo_monitor_1741;
    df_fifo_intf fifo_intf_1742(clock,reset);
    assign fifo_intf_1742.rd_en = AESL_inst_myproject.layer3_out_389_U.if_read & AESL_inst_myproject.layer3_out_389_U.if_empty_n;
    assign fifo_intf_1742.wr_en = AESL_inst_myproject.layer3_out_389_U.if_write & AESL_inst_myproject.layer3_out_389_U.if_full_n;
    assign fifo_intf_1742.fifo_rd_block = 0;
    assign fifo_intf_1742.fifo_wr_block = 0;
    assign fifo_intf_1742.finish = finish;
    csv_file_dump fifo_csv_dumper_1742;
    csv_file_dump cstatus_csv_dumper_1742;
    df_fifo_monitor fifo_monitor_1742;
    df_fifo_intf fifo_intf_1743(clock,reset);
    assign fifo_intf_1743.rd_en = AESL_inst_myproject.layer3_out_390_U.if_read & AESL_inst_myproject.layer3_out_390_U.if_empty_n;
    assign fifo_intf_1743.wr_en = AESL_inst_myproject.layer3_out_390_U.if_write & AESL_inst_myproject.layer3_out_390_U.if_full_n;
    assign fifo_intf_1743.fifo_rd_block = 0;
    assign fifo_intf_1743.fifo_wr_block = 0;
    assign fifo_intf_1743.finish = finish;
    csv_file_dump fifo_csv_dumper_1743;
    csv_file_dump cstatus_csv_dumper_1743;
    df_fifo_monitor fifo_monitor_1743;
    df_fifo_intf fifo_intf_1744(clock,reset);
    assign fifo_intf_1744.rd_en = AESL_inst_myproject.layer3_out_391_U.if_read & AESL_inst_myproject.layer3_out_391_U.if_empty_n;
    assign fifo_intf_1744.wr_en = AESL_inst_myproject.layer3_out_391_U.if_write & AESL_inst_myproject.layer3_out_391_U.if_full_n;
    assign fifo_intf_1744.fifo_rd_block = 0;
    assign fifo_intf_1744.fifo_wr_block = 0;
    assign fifo_intf_1744.finish = finish;
    csv_file_dump fifo_csv_dumper_1744;
    csv_file_dump cstatus_csv_dumper_1744;
    df_fifo_monitor fifo_monitor_1744;
    df_fifo_intf fifo_intf_1745(clock,reset);
    assign fifo_intf_1745.rd_en = AESL_inst_myproject.layer3_out_392_U.if_read & AESL_inst_myproject.layer3_out_392_U.if_empty_n;
    assign fifo_intf_1745.wr_en = AESL_inst_myproject.layer3_out_392_U.if_write & AESL_inst_myproject.layer3_out_392_U.if_full_n;
    assign fifo_intf_1745.fifo_rd_block = 0;
    assign fifo_intf_1745.fifo_wr_block = 0;
    assign fifo_intf_1745.finish = finish;
    csv_file_dump fifo_csv_dumper_1745;
    csv_file_dump cstatus_csv_dumper_1745;
    df_fifo_monitor fifo_monitor_1745;
    df_fifo_intf fifo_intf_1746(clock,reset);
    assign fifo_intf_1746.rd_en = AESL_inst_myproject.layer3_out_393_U.if_read & AESL_inst_myproject.layer3_out_393_U.if_empty_n;
    assign fifo_intf_1746.wr_en = AESL_inst_myproject.layer3_out_393_U.if_write & AESL_inst_myproject.layer3_out_393_U.if_full_n;
    assign fifo_intf_1746.fifo_rd_block = 0;
    assign fifo_intf_1746.fifo_wr_block = 0;
    assign fifo_intf_1746.finish = finish;
    csv_file_dump fifo_csv_dumper_1746;
    csv_file_dump cstatus_csv_dumper_1746;
    df_fifo_monitor fifo_monitor_1746;
    df_fifo_intf fifo_intf_1747(clock,reset);
    assign fifo_intf_1747.rd_en = AESL_inst_myproject.layer3_out_394_U.if_read & AESL_inst_myproject.layer3_out_394_U.if_empty_n;
    assign fifo_intf_1747.wr_en = AESL_inst_myproject.layer3_out_394_U.if_write & AESL_inst_myproject.layer3_out_394_U.if_full_n;
    assign fifo_intf_1747.fifo_rd_block = 0;
    assign fifo_intf_1747.fifo_wr_block = 0;
    assign fifo_intf_1747.finish = finish;
    csv_file_dump fifo_csv_dumper_1747;
    csv_file_dump cstatus_csv_dumper_1747;
    df_fifo_monitor fifo_monitor_1747;
    df_fifo_intf fifo_intf_1748(clock,reset);
    assign fifo_intf_1748.rd_en = AESL_inst_myproject.layer3_out_395_U.if_read & AESL_inst_myproject.layer3_out_395_U.if_empty_n;
    assign fifo_intf_1748.wr_en = AESL_inst_myproject.layer3_out_395_U.if_write & AESL_inst_myproject.layer3_out_395_U.if_full_n;
    assign fifo_intf_1748.fifo_rd_block = 0;
    assign fifo_intf_1748.fifo_wr_block = 0;
    assign fifo_intf_1748.finish = finish;
    csv_file_dump fifo_csv_dumper_1748;
    csv_file_dump cstatus_csv_dumper_1748;
    df_fifo_monitor fifo_monitor_1748;
    df_fifo_intf fifo_intf_1749(clock,reset);
    assign fifo_intf_1749.rd_en = AESL_inst_myproject.layer3_out_396_U.if_read & AESL_inst_myproject.layer3_out_396_U.if_empty_n;
    assign fifo_intf_1749.wr_en = AESL_inst_myproject.layer3_out_396_U.if_write & AESL_inst_myproject.layer3_out_396_U.if_full_n;
    assign fifo_intf_1749.fifo_rd_block = 0;
    assign fifo_intf_1749.fifo_wr_block = 0;
    assign fifo_intf_1749.finish = finish;
    csv_file_dump fifo_csv_dumper_1749;
    csv_file_dump cstatus_csv_dumper_1749;
    df_fifo_monitor fifo_monitor_1749;
    df_fifo_intf fifo_intf_1750(clock,reset);
    assign fifo_intf_1750.rd_en = AESL_inst_myproject.layer3_out_397_U.if_read & AESL_inst_myproject.layer3_out_397_U.if_empty_n;
    assign fifo_intf_1750.wr_en = AESL_inst_myproject.layer3_out_397_U.if_write & AESL_inst_myproject.layer3_out_397_U.if_full_n;
    assign fifo_intf_1750.fifo_rd_block = 0;
    assign fifo_intf_1750.fifo_wr_block = 0;
    assign fifo_intf_1750.finish = finish;
    csv_file_dump fifo_csv_dumper_1750;
    csv_file_dump cstatus_csv_dumper_1750;
    df_fifo_monitor fifo_monitor_1750;
    df_fifo_intf fifo_intf_1751(clock,reset);
    assign fifo_intf_1751.rd_en = AESL_inst_myproject.layer3_out_398_U.if_read & AESL_inst_myproject.layer3_out_398_U.if_empty_n;
    assign fifo_intf_1751.wr_en = AESL_inst_myproject.layer3_out_398_U.if_write & AESL_inst_myproject.layer3_out_398_U.if_full_n;
    assign fifo_intf_1751.fifo_rd_block = 0;
    assign fifo_intf_1751.fifo_wr_block = 0;
    assign fifo_intf_1751.finish = finish;
    csv_file_dump fifo_csv_dumper_1751;
    csv_file_dump cstatus_csv_dumper_1751;
    df_fifo_monitor fifo_monitor_1751;
    df_fifo_intf fifo_intf_1752(clock,reset);
    assign fifo_intf_1752.rd_en = AESL_inst_myproject.layer3_out_399_U.if_read & AESL_inst_myproject.layer3_out_399_U.if_empty_n;
    assign fifo_intf_1752.wr_en = AESL_inst_myproject.layer3_out_399_U.if_write & AESL_inst_myproject.layer3_out_399_U.if_full_n;
    assign fifo_intf_1752.fifo_rd_block = 0;
    assign fifo_intf_1752.fifo_wr_block = 0;
    assign fifo_intf_1752.finish = finish;
    csv_file_dump fifo_csv_dumper_1752;
    csv_file_dump cstatus_csv_dumper_1752;
    df_fifo_monitor fifo_monitor_1752;
    df_fifo_intf fifo_intf_1753(clock,reset);
    assign fifo_intf_1753.rd_en = AESL_inst_myproject.layer3_out_400_U.if_read & AESL_inst_myproject.layer3_out_400_U.if_empty_n;
    assign fifo_intf_1753.wr_en = AESL_inst_myproject.layer3_out_400_U.if_write & AESL_inst_myproject.layer3_out_400_U.if_full_n;
    assign fifo_intf_1753.fifo_rd_block = 0;
    assign fifo_intf_1753.fifo_wr_block = 0;
    assign fifo_intf_1753.finish = finish;
    csv_file_dump fifo_csv_dumper_1753;
    csv_file_dump cstatus_csv_dumper_1753;
    df_fifo_monitor fifo_monitor_1753;
    df_fifo_intf fifo_intf_1754(clock,reset);
    assign fifo_intf_1754.rd_en = AESL_inst_myproject.layer3_out_401_U.if_read & AESL_inst_myproject.layer3_out_401_U.if_empty_n;
    assign fifo_intf_1754.wr_en = AESL_inst_myproject.layer3_out_401_U.if_write & AESL_inst_myproject.layer3_out_401_U.if_full_n;
    assign fifo_intf_1754.fifo_rd_block = 0;
    assign fifo_intf_1754.fifo_wr_block = 0;
    assign fifo_intf_1754.finish = finish;
    csv_file_dump fifo_csv_dumper_1754;
    csv_file_dump cstatus_csv_dumper_1754;
    df_fifo_monitor fifo_monitor_1754;
    df_fifo_intf fifo_intf_1755(clock,reset);
    assign fifo_intf_1755.rd_en = AESL_inst_myproject.layer3_out_402_U.if_read & AESL_inst_myproject.layer3_out_402_U.if_empty_n;
    assign fifo_intf_1755.wr_en = AESL_inst_myproject.layer3_out_402_U.if_write & AESL_inst_myproject.layer3_out_402_U.if_full_n;
    assign fifo_intf_1755.fifo_rd_block = 0;
    assign fifo_intf_1755.fifo_wr_block = 0;
    assign fifo_intf_1755.finish = finish;
    csv_file_dump fifo_csv_dumper_1755;
    csv_file_dump cstatus_csv_dumper_1755;
    df_fifo_monitor fifo_monitor_1755;
    df_fifo_intf fifo_intf_1756(clock,reset);
    assign fifo_intf_1756.rd_en = AESL_inst_myproject.layer3_out_403_U.if_read & AESL_inst_myproject.layer3_out_403_U.if_empty_n;
    assign fifo_intf_1756.wr_en = AESL_inst_myproject.layer3_out_403_U.if_write & AESL_inst_myproject.layer3_out_403_U.if_full_n;
    assign fifo_intf_1756.fifo_rd_block = 0;
    assign fifo_intf_1756.fifo_wr_block = 0;
    assign fifo_intf_1756.finish = finish;
    csv_file_dump fifo_csv_dumper_1756;
    csv_file_dump cstatus_csv_dumper_1756;
    df_fifo_monitor fifo_monitor_1756;
    df_fifo_intf fifo_intf_1757(clock,reset);
    assign fifo_intf_1757.rd_en = AESL_inst_myproject.layer3_out_404_U.if_read & AESL_inst_myproject.layer3_out_404_U.if_empty_n;
    assign fifo_intf_1757.wr_en = AESL_inst_myproject.layer3_out_404_U.if_write & AESL_inst_myproject.layer3_out_404_U.if_full_n;
    assign fifo_intf_1757.fifo_rd_block = 0;
    assign fifo_intf_1757.fifo_wr_block = 0;
    assign fifo_intf_1757.finish = finish;
    csv_file_dump fifo_csv_dumper_1757;
    csv_file_dump cstatus_csv_dumper_1757;
    df_fifo_monitor fifo_monitor_1757;
    df_fifo_intf fifo_intf_1758(clock,reset);
    assign fifo_intf_1758.rd_en = AESL_inst_myproject.layer3_out_405_U.if_read & AESL_inst_myproject.layer3_out_405_U.if_empty_n;
    assign fifo_intf_1758.wr_en = AESL_inst_myproject.layer3_out_405_U.if_write & AESL_inst_myproject.layer3_out_405_U.if_full_n;
    assign fifo_intf_1758.fifo_rd_block = 0;
    assign fifo_intf_1758.fifo_wr_block = 0;
    assign fifo_intf_1758.finish = finish;
    csv_file_dump fifo_csv_dumper_1758;
    csv_file_dump cstatus_csv_dumper_1758;
    df_fifo_monitor fifo_monitor_1758;
    df_fifo_intf fifo_intf_1759(clock,reset);
    assign fifo_intf_1759.rd_en = AESL_inst_myproject.layer3_out_406_U.if_read & AESL_inst_myproject.layer3_out_406_U.if_empty_n;
    assign fifo_intf_1759.wr_en = AESL_inst_myproject.layer3_out_406_U.if_write & AESL_inst_myproject.layer3_out_406_U.if_full_n;
    assign fifo_intf_1759.fifo_rd_block = 0;
    assign fifo_intf_1759.fifo_wr_block = 0;
    assign fifo_intf_1759.finish = finish;
    csv_file_dump fifo_csv_dumper_1759;
    csv_file_dump cstatus_csv_dumper_1759;
    df_fifo_monitor fifo_monitor_1759;
    df_fifo_intf fifo_intf_1760(clock,reset);
    assign fifo_intf_1760.rd_en = AESL_inst_myproject.layer3_out_407_U.if_read & AESL_inst_myproject.layer3_out_407_U.if_empty_n;
    assign fifo_intf_1760.wr_en = AESL_inst_myproject.layer3_out_407_U.if_write & AESL_inst_myproject.layer3_out_407_U.if_full_n;
    assign fifo_intf_1760.fifo_rd_block = 0;
    assign fifo_intf_1760.fifo_wr_block = 0;
    assign fifo_intf_1760.finish = finish;
    csv_file_dump fifo_csv_dumper_1760;
    csv_file_dump cstatus_csv_dumper_1760;
    df_fifo_monitor fifo_monitor_1760;
    df_fifo_intf fifo_intf_1761(clock,reset);
    assign fifo_intf_1761.rd_en = AESL_inst_myproject.layer3_out_408_U.if_read & AESL_inst_myproject.layer3_out_408_U.if_empty_n;
    assign fifo_intf_1761.wr_en = AESL_inst_myproject.layer3_out_408_U.if_write & AESL_inst_myproject.layer3_out_408_U.if_full_n;
    assign fifo_intf_1761.fifo_rd_block = 0;
    assign fifo_intf_1761.fifo_wr_block = 0;
    assign fifo_intf_1761.finish = finish;
    csv_file_dump fifo_csv_dumper_1761;
    csv_file_dump cstatus_csv_dumper_1761;
    df_fifo_monitor fifo_monitor_1761;
    df_fifo_intf fifo_intf_1762(clock,reset);
    assign fifo_intf_1762.rd_en = AESL_inst_myproject.layer3_out_409_U.if_read & AESL_inst_myproject.layer3_out_409_U.if_empty_n;
    assign fifo_intf_1762.wr_en = AESL_inst_myproject.layer3_out_409_U.if_write & AESL_inst_myproject.layer3_out_409_U.if_full_n;
    assign fifo_intf_1762.fifo_rd_block = 0;
    assign fifo_intf_1762.fifo_wr_block = 0;
    assign fifo_intf_1762.finish = finish;
    csv_file_dump fifo_csv_dumper_1762;
    csv_file_dump cstatus_csv_dumper_1762;
    df_fifo_monitor fifo_monitor_1762;
    df_fifo_intf fifo_intf_1763(clock,reset);
    assign fifo_intf_1763.rd_en = AESL_inst_myproject.layer3_out_410_U.if_read & AESL_inst_myproject.layer3_out_410_U.if_empty_n;
    assign fifo_intf_1763.wr_en = AESL_inst_myproject.layer3_out_410_U.if_write & AESL_inst_myproject.layer3_out_410_U.if_full_n;
    assign fifo_intf_1763.fifo_rd_block = 0;
    assign fifo_intf_1763.fifo_wr_block = 0;
    assign fifo_intf_1763.finish = finish;
    csv_file_dump fifo_csv_dumper_1763;
    csv_file_dump cstatus_csv_dumper_1763;
    df_fifo_monitor fifo_monitor_1763;
    df_fifo_intf fifo_intf_1764(clock,reset);
    assign fifo_intf_1764.rd_en = AESL_inst_myproject.layer3_out_411_U.if_read & AESL_inst_myproject.layer3_out_411_U.if_empty_n;
    assign fifo_intf_1764.wr_en = AESL_inst_myproject.layer3_out_411_U.if_write & AESL_inst_myproject.layer3_out_411_U.if_full_n;
    assign fifo_intf_1764.fifo_rd_block = 0;
    assign fifo_intf_1764.fifo_wr_block = 0;
    assign fifo_intf_1764.finish = finish;
    csv_file_dump fifo_csv_dumper_1764;
    csv_file_dump cstatus_csv_dumper_1764;
    df_fifo_monitor fifo_monitor_1764;
    df_fifo_intf fifo_intf_1765(clock,reset);
    assign fifo_intf_1765.rd_en = AESL_inst_myproject.layer3_out_412_U.if_read & AESL_inst_myproject.layer3_out_412_U.if_empty_n;
    assign fifo_intf_1765.wr_en = AESL_inst_myproject.layer3_out_412_U.if_write & AESL_inst_myproject.layer3_out_412_U.if_full_n;
    assign fifo_intf_1765.fifo_rd_block = 0;
    assign fifo_intf_1765.fifo_wr_block = 0;
    assign fifo_intf_1765.finish = finish;
    csv_file_dump fifo_csv_dumper_1765;
    csv_file_dump cstatus_csv_dumper_1765;
    df_fifo_monitor fifo_monitor_1765;
    df_fifo_intf fifo_intf_1766(clock,reset);
    assign fifo_intf_1766.rd_en = AESL_inst_myproject.layer3_out_413_U.if_read & AESL_inst_myproject.layer3_out_413_U.if_empty_n;
    assign fifo_intf_1766.wr_en = AESL_inst_myproject.layer3_out_413_U.if_write & AESL_inst_myproject.layer3_out_413_U.if_full_n;
    assign fifo_intf_1766.fifo_rd_block = 0;
    assign fifo_intf_1766.fifo_wr_block = 0;
    assign fifo_intf_1766.finish = finish;
    csv_file_dump fifo_csv_dumper_1766;
    csv_file_dump cstatus_csv_dumper_1766;
    df_fifo_monitor fifo_monitor_1766;
    df_fifo_intf fifo_intf_1767(clock,reset);
    assign fifo_intf_1767.rd_en = AESL_inst_myproject.layer3_out_414_U.if_read & AESL_inst_myproject.layer3_out_414_U.if_empty_n;
    assign fifo_intf_1767.wr_en = AESL_inst_myproject.layer3_out_414_U.if_write & AESL_inst_myproject.layer3_out_414_U.if_full_n;
    assign fifo_intf_1767.fifo_rd_block = 0;
    assign fifo_intf_1767.fifo_wr_block = 0;
    assign fifo_intf_1767.finish = finish;
    csv_file_dump fifo_csv_dumper_1767;
    csv_file_dump cstatus_csv_dumper_1767;
    df_fifo_monitor fifo_monitor_1767;
    df_fifo_intf fifo_intf_1768(clock,reset);
    assign fifo_intf_1768.rd_en = AESL_inst_myproject.layer3_out_415_U.if_read & AESL_inst_myproject.layer3_out_415_U.if_empty_n;
    assign fifo_intf_1768.wr_en = AESL_inst_myproject.layer3_out_415_U.if_write & AESL_inst_myproject.layer3_out_415_U.if_full_n;
    assign fifo_intf_1768.fifo_rd_block = 0;
    assign fifo_intf_1768.fifo_wr_block = 0;
    assign fifo_intf_1768.finish = finish;
    csv_file_dump fifo_csv_dumper_1768;
    csv_file_dump cstatus_csv_dumper_1768;
    df_fifo_monitor fifo_monitor_1768;
    df_fifo_intf fifo_intf_1769(clock,reset);
    assign fifo_intf_1769.rd_en = AESL_inst_myproject.layer3_out_416_U.if_read & AESL_inst_myproject.layer3_out_416_U.if_empty_n;
    assign fifo_intf_1769.wr_en = AESL_inst_myproject.layer3_out_416_U.if_write & AESL_inst_myproject.layer3_out_416_U.if_full_n;
    assign fifo_intf_1769.fifo_rd_block = 0;
    assign fifo_intf_1769.fifo_wr_block = 0;
    assign fifo_intf_1769.finish = finish;
    csv_file_dump fifo_csv_dumper_1769;
    csv_file_dump cstatus_csv_dumper_1769;
    df_fifo_monitor fifo_monitor_1769;
    df_fifo_intf fifo_intf_1770(clock,reset);
    assign fifo_intf_1770.rd_en = AESL_inst_myproject.layer3_out_417_U.if_read & AESL_inst_myproject.layer3_out_417_U.if_empty_n;
    assign fifo_intf_1770.wr_en = AESL_inst_myproject.layer3_out_417_U.if_write & AESL_inst_myproject.layer3_out_417_U.if_full_n;
    assign fifo_intf_1770.fifo_rd_block = 0;
    assign fifo_intf_1770.fifo_wr_block = 0;
    assign fifo_intf_1770.finish = finish;
    csv_file_dump fifo_csv_dumper_1770;
    csv_file_dump cstatus_csv_dumper_1770;
    df_fifo_monitor fifo_monitor_1770;
    df_fifo_intf fifo_intf_1771(clock,reset);
    assign fifo_intf_1771.rd_en = AESL_inst_myproject.layer3_out_418_U.if_read & AESL_inst_myproject.layer3_out_418_U.if_empty_n;
    assign fifo_intf_1771.wr_en = AESL_inst_myproject.layer3_out_418_U.if_write & AESL_inst_myproject.layer3_out_418_U.if_full_n;
    assign fifo_intf_1771.fifo_rd_block = 0;
    assign fifo_intf_1771.fifo_wr_block = 0;
    assign fifo_intf_1771.finish = finish;
    csv_file_dump fifo_csv_dumper_1771;
    csv_file_dump cstatus_csv_dumper_1771;
    df_fifo_monitor fifo_monitor_1771;
    df_fifo_intf fifo_intf_1772(clock,reset);
    assign fifo_intf_1772.rd_en = AESL_inst_myproject.layer3_out_419_U.if_read & AESL_inst_myproject.layer3_out_419_U.if_empty_n;
    assign fifo_intf_1772.wr_en = AESL_inst_myproject.layer3_out_419_U.if_write & AESL_inst_myproject.layer3_out_419_U.if_full_n;
    assign fifo_intf_1772.fifo_rd_block = 0;
    assign fifo_intf_1772.fifo_wr_block = 0;
    assign fifo_intf_1772.finish = finish;
    csv_file_dump fifo_csv_dumper_1772;
    csv_file_dump cstatus_csv_dumper_1772;
    df_fifo_monitor fifo_monitor_1772;
    df_fifo_intf fifo_intf_1773(clock,reset);
    assign fifo_intf_1773.rd_en = AESL_inst_myproject.layer3_out_420_U.if_read & AESL_inst_myproject.layer3_out_420_U.if_empty_n;
    assign fifo_intf_1773.wr_en = AESL_inst_myproject.layer3_out_420_U.if_write & AESL_inst_myproject.layer3_out_420_U.if_full_n;
    assign fifo_intf_1773.fifo_rd_block = 0;
    assign fifo_intf_1773.fifo_wr_block = 0;
    assign fifo_intf_1773.finish = finish;
    csv_file_dump fifo_csv_dumper_1773;
    csv_file_dump cstatus_csv_dumper_1773;
    df_fifo_monitor fifo_monitor_1773;
    df_fifo_intf fifo_intf_1774(clock,reset);
    assign fifo_intf_1774.rd_en = AESL_inst_myproject.layer3_out_421_U.if_read & AESL_inst_myproject.layer3_out_421_U.if_empty_n;
    assign fifo_intf_1774.wr_en = AESL_inst_myproject.layer3_out_421_U.if_write & AESL_inst_myproject.layer3_out_421_U.if_full_n;
    assign fifo_intf_1774.fifo_rd_block = 0;
    assign fifo_intf_1774.fifo_wr_block = 0;
    assign fifo_intf_1774.finish = finish;
    csv_file_dump fifo_csv_dumper_1774;
    csv_file_dump cstatus_csv_dumper_1774;
    df_fifo_monitor fifo_monitor_1774;
    df_fifo_intf fifo_intf_1775(clock,reset);
    assign fifo_intf_1775.rd_en = AESL_inst_myproject.layer3_out_422_U.if_read & AESL_inst_myproject.layer3_out_422_U.if_empty_n;
    assign fifo_intf_1775.wr_en = AESL_inst_myproject.layer3_out_422_U.if_write & AESL_inst_myproject.layer3_out_422_U.if_full_n;
    assign fifo_intf_1775.fifo_rd_block = 0;
    assign fifo_intf_1775.fifo_wr_block = 0;
    assign fifo_intf_1775.finish = finish;
    csv_file_dump fifo_csv_dumper_1775;
    csv_file_dump cstatus_csv_dumper_1775;
    df_fifo_monitor fifo_monitor_1775;
    df_fifo_intf fifo_intf_1776(clock,reset);
    assign fifo_intf_1776.rd_en = AESL_inst_myproject.layer3_out_423_U.if_read & AESL_inst_myproject.layer3_out_423_U.if_empty_n;
    assign fifo_intf_1776.wr_en = AESL_inst_myproject.layer3_out_423_U.if_write & AESL_inst_myproject.layer3_out_423_U.if_full_n;
    assign fifo_intf_1776.fifo_rd_block = 0;
    assign fifo_intf_1776.fifo_wr_block = 0;
    assign fifo_intf_1776.finish = finish;
    csv_file_dump fifo_csv_dumper_1776;
    csv_file_dump cstatus_csv_dumper_1776;
    df_fifo_monitor fifo_monitor_1776;
    df_fifo_intf fifo_intf_1777(clock,reset);
    assign fifo_intf_1777.rd_en = AESL_inst_myproject.layer3_out_424_U.if_read & AESL_inst_myproject.layer3_out_424_U.if_empty_n;
    assign fifo_intf_1777.wr_en = AESL_inst_myproject.layer3_out_424_U.if_write & AESL_inst_myproject.layer3_out_424_U.if_full_n;
    assign fifo_intf_1777.fifo_rd_block = 0;
    assign fifo_intf_1777.fifo_wr_block = 0;
    assign fifo_intf_1777.finish = finish;
    csv_file_dump fifo_csv_dumper_1777;
    csv_file_dump cstatus_csv_dumper_1777;
    df_fifo_monitor fifo_monitor_1777;
    df_fifo_intf fifo_intf_1778(clock,reset);
    assign fifo_intf_1778.rd_en = AESL_inst_myproject.layer3_out_425_U.if_read & AESL_inst_myproject.layer3_out_425_U.if_empty_n;
    assign fifo_intf_1778.wr_en = AESL_inst_myproject.layer3_out_425_U.if_write & AESL_inst_myproject.layer3_out_425_U.if_full_n;
    assign fifo_intf_1778.fifo_rd_block = 0;
    assign fifo_intf_1778.fifo_wr_block = 0;
    assign fifo_intf_1778.finish = finish;
    csv_file_dump fifo_csv_dumper_1778;
    csv_file_dump cstatus_csv_dumper_1778;
    df_fifo_monitor fifo_monitor_1778;
    df_fifo_intf fifo_intf_1779(clock,reset);
    assign fifo_intf_1779.rd_en = AESL_inst_myproject.layer3_out_426_U.if_read & AESL_inst_myproject.layer3_out_426_U.if_empty_n;
    assign fifo_intf_1779.wr_en = AESL_inst_myproject.layer3_out_426_U.if_write & AESL_inst_myproject.layer3_out_426_U.if_full_n;
    assign fifo_intf_1779.fifo_rd_block = 0;
    assign fifo_intf_1779.fifo_wr_block = 0;
    assign fifo_intf_1779.finish = finish;
    csv_file_dump fifo_csv_dumper_1779;
    csv_file_dump cstatus_csv_dumper_1779;
    df_fifo_monitor fifo_monitor_1779;
    df_fifo_intf fifo_intf_1780(clock,reset);
    assign fifo_intf_1780.rd_en = AESL_inst_myproject.layer3_out_427_U.if_read & AESL_inst_myproject.layer3_out_427_U.if_empty_n;
    assign fifo_intf_1780.wr_en = AESL_inst_myproject.layer3_out_427_U.if_write & AESL_inst_myproject.layer3_out_427_U.if_full_n;
    assign fifo_intf_1780.fifo_rd_block = 0;
    assign fifo_intf_1780.fifo_wr_block = 0;
    assign fifo_intf_1780.finish = finish;
    csv_file_dump fifo_csv_dumper_1780;
    csv_file_dump cstatus_csv_dumper_1780;
    df_fifo_monitor fifo_monitor_1780;
    df_fifo_intf fifo_intf_1781(clock,reset);
    assign fifo_intf_1781.rd_en = AESL_inst_myproject.layer3_out_428_U.if_read & AESL_inst_myproject.layer3_out_428_U.if_empty_n;
    assign fifo_intf_1781.wr_en = AESL_inst_myproject.layer3_out_428_U.if_write & AESL_inst_myproject.layer3_out_428_U.if_full_n;
    assign fifo_intf_1781.fifo_rd_block = 0;
    assign fifo_intf_1781.fifo_wr_block = 0;
    assign fifo_intf_1781.finish = finish;
    csv_file_dump fifo_csv_dumper_1781;
    csv_file_dump cstatus_csv_dumper_1781;
    df_fifo_monitor fifo_monitor_1781;
    df_fifo_intf fifo_intf_1782(clock,reset);
    assign fifo_intf_1782.rd_en = AESL_inst_myproject.layer3_out_429_U.if_read & AESL_inst_myproject.layer3_out_429_U.if_empty_n;
    assign fifo_intf_1782.wr_en = AESL_inst_myproject.layer3_out_429_U.if_write & AESL_inst_myproject.layer3_out_429_U.if_full_n;
    assign fifo_intf_1782.fifo_rd_block = 0;
    assign fifo_intf_1782.fifo_wr_block = 0;
    assign fifo_intf_1782.finish = finish;
    csv_file_dump fifo_csv_dumper_1782;
    csv_file_dump cstatus_csv_dumper_1782;
    df_fifo_monitor fifo_monitor_1782;
    df_fifo_intf fifo_intf_1783(clock,reset);
    assign fifo_intf_1783.rd_en = AESL_inst_myproject.layer3_out_430_U.if_read & AESL_inst_myproject.layer3_out_430_U.if_empty_n;
    assign fifo_intf_1783.wr_en = AESL_inst_myproject.layer3_out_430_U.if_write & AESL_inst_myproject.layer3_out_430_U.if_full_n;
    assign fifo_intf_1783.fifo_rd_block = 0;
    assign fifo_intf_1783.fifo_wr_block = 0;
    assign fifo_intf_1783.finish = finish;
    csv_file_dump fifo_csv_dumper_1783;
    csv_file_dump cstatus_csv_dumper_1783;
    df_fifo_monitor fifo_monitor_1783;
    df_fifo_intf fifo_intf_1784(clock,reset);
    assign fifo_intf_1784.rd_en = AESL_inst_myproject.layer3_out_431_U.if_read & AESL_inst_myproject.layer3_out_431_U.if_empty_n;
    assign fifo_intf_1784.wr_en = AESL_inst_myproject.layer3_out_431_U.if_write & AESL_inst_myproject.layer3_out_431_U.if_full_n;
    assign fifo_intf_1784.fifo_rd_block = 0;
    assign fifo_intf_1784.fifo_wr_block = 0;
    assign fifo_intf_1784.finish = finish;
    csv_file_dump fifo_csv_dumper_1784;
    csv_file_dump cstatus_csv_dumper_1784;
    df_fifo_monitor fifo_monitor_1784;
    df_fifo_intf fifo_intf_1785(clock,reset);
    assign fifo_intf_1785.rd_en = AESL_inst_myproject.layer3_out_432_U.if_read & AESL_inst_myproject.layer3_out_432_U.if_empty_n;
    assign fifo_intf_1785.wr_en = AESL_inst_myproject.layer3_out_432_U.if_write & AESL_inst_myproject.layer3_out_432_U.if_full_n;
    assign fifo_intf_1785.fifo_rd_block = 0;
    assign fifo_intf_1785.fifo_wr_block = 0;
    assign fifo_intf_1785.finish = finish;
    csv_file_dump fifo_csv_dumper_1785;
    csv_file_dump cstatus_csv_dumper_1785;
    df_fifo_monitor fifo_monitor_1785;
    df_fifo_intf fifo_intf_1786(clock,reset);
    assign fifo_intf_1786.rd_en = AESL_inst_myproject.layer3_out_433_U.if_read & AESL_inst_myproject.layer3_out_433_U.if_empty_n;
    assign fifo_intf_1786.wr_en = AESL_inst_myproject.layer3_out_433_U.if_write & AESL_inst_myproject.layer3_out_433_U.if_full_n;
    assign fifo_intf_1786.fifo_rd_block = 0;
    assign fifo_intf_1786.fifo_wr_block = 0;
    assign fifo_intf_1786.finish = finish;
    csv_file_dump fifo_csv_dumper_1786;
    csv_file_dump cstatus_csv_dumper_1786;
    df_fifo_monitor fifo_monitor_1786;
    df_fifo_intf fifo_intf_1787(clock,reset);
    assign fifo_intf_1787.rd_en = AESL_inst_myproject.layer3_out_434_U.if_read & AESL_inst_myproject.layer3_out_434_U.if_empty_n;
    assign fifo_intf_1787.wr_en = AESL_inst_myproject.layer3_out_434_U.if_write & AESL_inst_myproject.layer3_out_434_U.if_full_n;
    assign fifo_intf_1787.fifo_rd_block = 0;
    assign fifo_intf_1787.fifo_wr_block = 0;
    assign fifo_intf_1787.finish = finish;
    csv_file_dump fifo_csv_dumper_1787;
    csv_file_dump cstatus_csv_dumper_1787;
    df_fifo_monitor fifo_monitor_1787;
    df_fifo_intf fifo_intf_1788(clock,reset);
    assign fifo_intf_1788.rd_en = AESL_inst_myproject.layer3_out_435_U.if_read & AESL_inst_myproject.layer3_out_435_U.if_empty_n;
    assign fifo_intf_1788.wr_en = AESL_inst_myproject.layer3_out_435_U.if_write & AESL_inst_myproject.layer3_out_435_U.if_full_n;
    assign fifo_intf_1788.fifo_rd_block = 0;
    assign fifo_intf_1788.fifo_wr_block = 0;
    assign fifo_intf_1788.finish = finish;
    csv_file_dump fifo_csv_dumper_1788;
    csv_file_dump cstatus_csv_dumper_1788;
    df_fifo_monitor fifo_monitor_1788;
    df_fifo_intf fifo_intf_1789(clock,reset);
    assign fifo_intf_1789.rd_en = AESL_inst_myproject.layer3_out_436_U.if_read & AESL_inst_myproject.layer3_out_436_U.if_empty_n;
    assign fifo_intf_1789.wr_en = AESL_inst_myproject.layer3_out_436_U.if_write & AESL_inst_myproject.layer3_out_436_U.if_full_n;
    assign fifo_intf_1789.fifo_rd_block = 0;
    assign fifo_intf_1789.fifo_wr_block = 0;
    assign fifo_intf_1789.finish = finish;
    csv_file_dump fifo_csv_dumper_1789;
    csv_file_dump cstatus_csv_dumper_1789;
    df_fifo_monitor fifo_monitor_1789;
    df_fifo_intf fifo_intf_1790(clock,reset);
    assign fifo_intf_1790.rd_en = AESL_inst_myproject.layer3_out_437_U.if_read & AESL_inst_myproject.layer3_out_437_U.if_empty_n;
    assign fifo_intf_1790.wr_en = AESL_inst_myproject.layer3_out_437_U.if_write & AESL_inst_myproject.layer3_out_437_U.if_full_n;
    assign fifo_intf_1790.fifo_rd_block = 0;
    assign fifo_intf_1790.fifo_wr_block = 0;
    assign fifo_intf_1790.finish = finish;
    csv_file_dump fifo_csv_dumper_1790;
    csv_file_dump cstatus_csv_dumper_1790;
    df_fifo_monitor fifo_monitor_1790;
    df_fifo_intf fifo_intf_1791(clock,reset);
    assign fifo_intf_1791.rd_en = AESL_inst_myproject.layer3_out_438_U.if_read & AESL_inst_myproject.layer3_out_438_U.if_empty_n;
    assign fifo_intf_1791.wr_en = AESL_inst_myproject.layer3_out_438_U.if_write & AESL_inst_myproject.layer3_out_438_U.if_full_n;
    assign fifo_intf_1791.fifo_rd_block = 0;
    assign fifo_intf_1791.fifo_wr_block = 0;
    assign fifo_intf_1791.finish = finish;
    csv_file_dump fifo_csv_dumper_1791;
    csv_file_dump cstatus_csv_dumper_1791;
    df_fifo_monitor fifo_monitor_1791;
    df_fifo_intf fifo_intf_1792(clock,reset);
    assign fifo_intf_1792.rd_en = AESL_inst_myproject.layer3_out_439_U.if_read & AESL_inst_myproject.layer3_out_439_U.if_empty_n;
    assign fifo_intf_1792.wr_en = AESL_inst_myproject.layer3_out_439_U.if_write & AESL_inst_myproject.layer3_out_439_U.if_full_n;
    assign fifo_intf_1792.fifo_rd_block = 0;
    assign fifo_intf_1792.fifo_wr_block = 0;
    assign fifo_intf_1792.finish = finish;
    csv_file_dump fifo_csv_dumper_1792;
    csv_file_dump cstatus_csv_dumper_1792;
    df_fifo_monitor fifo_monitor_1792;
    df_fifo_intf fifo_intf_1793(clock,reset);
    assign fifo_intf_1793.rd_en = AESL_inst_myproject.layer3_out_440_U.if_read & AESL_inst_myproject.layer3_out_440_U.if_empty_n;
    assign fifo_intf_1793.wr_en = AESL_inst_myproject.layer3_out_440_U.if_write & AESL_inst_myproject.layer3_out_440_U.if_full_n;
    assign fifo_intf_1793.fifo_rd_block = 0;
    assign fifo_intf_1793.fifo_wr_block = 0;
    assign fifo_intf_1793.finish = finish;
    csv_file_dump fifo_csv_dumper_1793;
    csv_file_dump cstatus_csv_dumper_1793;
    df_fifo_monitor fifo_monitor_1793;
    df_fifo_intf fifo_intf_1794(clock,reset);
    assign fifo_intf_1794.rd_en = AESL_inst_myproject.layer3_out_441_U.if_read & AESL_inst_myproject.layer3_out_441_U.if_empty_n;
    assign fifo_intf_1794.wr_en = AESL_inst_myproject.layer3_out_441_U.if_write & AESL_inst_myproject.layer3_out_441_U.if_full_n;
    assign fifo_intf_1794.fifo_rd_block = 0;
    assign fifo_intf_1794.fifo_wr_block = 0;
    assign fifo_intf_1794.finish = finish;
    csv_file_dump fifo_csv_dumper_1794;
    csv_file_dump cstatus_csv_dumper_1794;
    df_fifo_monitor fifo_monitor_1794;
    df_fifo_intf fifo_intf_1795(clock,reset);
    assign fifo_intf_1795.rd_en = AESL_inst_myproject.layer3_out_442_U.if_read & AESL_inst_myproject.layer3_out_442_U.if_empty_n;
    assign fifo_intf_1795.wr_en = AESL_inst_myproject.layer3_out_442_U.if_write & AESL_inst_myproject.layer3_out_442_U.if_full_n;
    assign fifo_intf_1795.fifo_rd_block = 0;
    assign fifo_intf_1795.fifo_wr_block = 0;
    assign fifo_intf_1795.finish = finish;
    csv_file_dump fifo_csv_dumper_1795;
    csv_file_dump cstatus_csv_dumper_1795;
    df_fifo_monitor fifo_monitor_1795;
    df_fifo_intf fifo_intf_1796(clock,reset);
    assign fifo_intf_1796.rd_en = AESL_inst_myproject.layer3_out_443_U.if_read & AESL_inst_myproject.layer3_out_443_U.if_empty_n;
    assign fifo_intf_1796.wr_en = AESL_inst_myproject.layer3_out_443_U.if_write & AESL_inst_myproject.layer3_out_443_U.if_full_n;
    assign fifo_intf_1796.fifo_rd_block = 0;
    assign fifo_intf_1796.fifo_wr_block = 0;
    assign fifo_intf_1796.finish = finish;
    csv_file_dump fifo_csv_dumper_1796;
    csv_file_dump cstatus_csv_dumper_1796;
    df_fifo_monitor fifo_monitor_1796;
    df_fifo_intf fifo_intf_1797(clock,reset);
    assign fifo_intf_1797.rd_en = AESL_inst_myproject.layer3_out_444_U.if_read & AESL_inst_myproject.layer3_out_444_U.if_empty_n;
    assign fifo_intf_1797.wr_en = AESL_inst_myproject.layer3_out_444_U.if_write & AESL_inst_myproject.layer3_out_444_U.if_full_n;
    assign fifo_intf_1797.fifo_rd_block = 0;
    assign fifo_intf_1797.fifo_wr_block = 0;
    assign fifo_intf_1797.finish = finish;
    csv_file_dump fifo_csv_dumper_1797;
    csv_file_dump cstatus_csv_dumper_1797;
    df_fifo_monitor fifo_monitor_1797;
    df_fifo_intf fifo_intf_1798(clock,reset);
    assign fifo_intf_1798.rd_en = AESL_inst_myproject.layer3_out_445_U.if_read & AESL_inst_myproject.layer3_out_445_U.if_empty_n;
    assign fifo_intf_1798.wr_en = AESL_inst_myproject.layer3_out_445_U.if_write & AESL_inst_myproject.layer3_out_445_U.if_full_n;
    assign fifo_intf_1798.fifo_rd_block = 0;
    assign fifo_intf_1798.fifo_wr_block = 0;
    assign fifo_intf_1798.finish = finish;
    csv_file_dump fifo_csv_dumper_1798;
    csv_file_dump cstatus_csv_dumper_1798;
    df_fifo_monitor fifo_monitor_1798;
    df_fifo_intf fifo_intf_1799(clock,reset);
    assign fifo_intf_1799.rd_en = AESL_inst_myproject.layer3_out_446_U.if_read & AESL_inst_myproject.layer3_out_446_U.if_empty_n;
    assign fifo_intf_1799.wr_en = AESL_inst_myproject.layer3_out_446_U.if_write & AESL_inst_myproject.layer3_out_446_U.if_full_n;
    assign fifo_intf_1799.fifo_rd_block = 0;
    assign fifo_intf_1799.fifo_wr_block = 0;
    assign fifo_intf_1799.finish = finish;
    csv_file_dump fifo_csv_dumper_1799;
    csv_file_dump cstatus_csv_dumper_1799;
    df_fifo_monitor fifo_monitor_1799;
    df_fifo_intf fifo_intf_1800(clock,reset);
    assign fifo_intf_1800.rd_en = AESL_inst_myproject.layer3_out_447_U.if_read & AESL_inst_myproject.layer3_out_447_U.if_empty_n;
    assign fifo_intf_1800.wr_en = AESL_inst_myproject.layer3_out_447_U.if_write & AESL_inst_myproject.layer3_out_447_U.if_full_n;
    assign fifo_intf_1800.fifo_rd_block = 0;
    assign fifo_intf_1800.fifo_wr_block = 0;
    assign fifo_intf_1800.finish = finish;
    csv_file_dump fifo_csv_dumper_1800;
    csv_file_dump cstatus_csv_dumper_1800;
    df_fifo_monitor fifo_monitor_1800;
    df_fifo_intf fifo_intf_1801(clock,reset);
    assign fifo_intf_1801.rd_en = AESL_inst_myproject.layer3_out_448_U.if_read & AESL_inst_myproject.layer3_out_448_U.if_empty_n;
    assign fifo_intf_1801.wr_en = AESL_inst_myproject.layer3_out_448_U.if_write & AESL_inst_myproject.layer3_out_448_U.if_full_n;
    assign fifo_intf_1801.fifo_rd_block = 0;
    assign fifo_intf_1801.fifo_wr_block = 0;
    assign fifo_intf_1801.finish = finish;
    csv_file_dump fifo_csv_dumper_1801;
    csv_file_dump cstatus_csv_dumper_1801;
    df_fifo_monitor fifo_monitor_1801;
    df_fifo_intf fifo_intf_1802(clock,reset);
    assign fifo_intf_1802.rd_en = AESL_inst_myproject.layer3_out_449_U.if_read & AESL_inst_myproject.layer3_out_449_U.if_empty_n;
    assign fifo_intf_1802.wr_en = AESL_inst_myproject.layer3_out_449_U.if_write & AESL_inst_myproject.layer3_out_449_U.if_full_n;
    assign fifo_intf_1802.fifo_rd_block = 0;
    assign fifo_intf_1802.fifo_wr_block = 0;
    assign fifo_intf_1802.finish = finish;
    csv_file_dump fifo_csv_dumper_1802;
    csv_file_dump cstatus_csv_dumper_1802;
    df_fifo_monitor fifo_monitor_1802;
    df_fifo_intf fifo_intf_1803(clock,reset);
    assign fifo_intf_1803.rd_en = AESL_inst_myproject.layer3_out_450_U.if_read & AESL_inst_myproject.layer3_out_450_U.if_empty_n;
    assign fifo_intf_1803.wr_en = AESL_inst_myproject.layer3_out_450_U.if_write & AESL_inst_myproject.layer3_out_450_U.if_full_n;
    assign fifo_intf_1803.fifo_rd_block = 0;
    assign fifo_intf_1803.fifo_wr_block = 0;
    assign fifo_intf_1803.finish = finish;
    csv_file_dump fifo_csv_dumper_1803;
    csv_file_dump cstatus_csv_dumper_1803;
    df_fifo_monitor fifo_monitor_1803;
    df_fifo_intf fifo_intf_1804(clock,reset);
    assign fifo_intf_1804.rd_en = AESL_inst_myproject.layer3_out_451_U.if_read & AESL_inst_myproject.layer3_out_451_U.if_empty_n;
    assign fifo_intf_1804.wr_en = AESL_inst_myproject.layer3_out_451_U.if_write & AESL_inst_myproject.layer3_out_451_U.if_full_n;
    assign fifo_intf_1804.fifo_rd_block = 0;
    assign fifo_intf_1804.fifo_wr_block = 0;
    assign fifo_intf_1804.finish = finish;
    csv_file_dump fifo_csv_dumper_1804;
    csv_file_dump cstatus_csv_dumper_1804;
    df_fifo_monitor fifo_monitor_1804;
    df_fifo_intf fifo_intf_1805(clock,reset);
    assign fifo_intf_1805.rd_en = AESL_inst_myproject.layer3_out_452_U.if_read & AESL_inst_myproject.layer3_out_452_U.if_empty_n;
    assign fifo_intf_1805.wr_en = AESL_inst_myproject.layer3_out_452_U.if_write & AESL_inst_myproject.layer3_out_452_U.if_full_n;
    assign fifo_intf_1805.fifo_rd_block = 0;
    assign fifo_intf_1805.fifo_wr_block = 0;
    assign fifo_intf_1805.finish = finish;
    csv_file_dump fifo_csv_dumper_1805;
    csv_file_dump cstatus_csv_dumper_1805;
    df_fifo_monitor fifo_monitor_1805;
    df_fifo_intf fifo_intf_1806(clock,reset);
    assign fifo_intf_1806.rd_en = AESL_inst_myproject.layer3_out_453_U.if_read & AESL_inst_myproject.layer3_out_453_U.if_empty_n;
    assign fifo_intf_1806.wr_en = AESL_inst_myproject.layer3_out_453_U.if_write & AESL_inst_myproject.layer3_out_453_U.if_full_n;
    assign fifo_intf_1806.fifo_rd_block = 0;
    assign fifo_intf_1806.fifo_wr_block = 0;
    assign fifo_intf_1806.finish = finish;
    csv_file_dump fifo_csv_dumper_1806;
    csv_file_dump cstatus_csv_dumper_1806;
    df_fifo_monitor fifo_monitor_1806;
    df_fifo_intf fifo_intf_1807(clock,reset);
    assign fifo_intf_1807.rd_en = AESL_inst_myproject.layer3_out_454_U.if_read & AESL_inst_myproject.layer3_out_454_U.if_empty_n;
    assign fifo_intf_1807.wr_en = AESL_inst_myproject.layer3_out_454_U.if_write & AESL_inst_myproject.layer3_out_454_U.if_full_n;
    assign fifo_intf_1807.fifo_rd_block = 0;
    assign fifo_intf_1807.fifo_wr_block = 0;
    assign fifo_intf_1807.finish = finish;
    csv_file_dump fifo_csv_dumper_1807;
    csv_file_dump cstatus_csv_dumper_1807;
    df_fifo_monitor fifo_monitor_1807;
    df_fifo_intf fifo_intf_1808(clock,reset);
    assign fifo_intf_1808.rd_en = AESL_inst_myproject.layer3_out_455_U.if_read & AESL_inst_myproject.layer3_out_455_U.if_empty_n;
    assign fifo_intf_1808.wr_en = AESL_inst_myproject.layer3_out_455_U.if_write & AESL_inst_myproject.layer3_out_455_U.if_full_n;
    assign fifo_intf_1808.fifo_rd_block = 0;
    assign fifo_intf_1808.fifo_wr_block = 0;
    assign fifo_intf_1808.finish = finish;
    csv_file_dump fifo_csv_dumper_1808;
    csv_file_dump cstatus_csv_dumper_1808;
    df_fifo_monitor fifo_monitor_1808;
    df_fifo_intf fifo_intf_1809(clock,reset);
    assign fifo_intf_1809.rd_en = AESL_inst_myproject.layer3_out_456_U.if_read & AESL_inst_myproject.layer3_out_456_U.if_empty_n;
    assign fifo_intf_1809.wr_en = AESL_inst_myproject.layer3_out_456_U.if_write & AESL_inst_myproject.layer3_out_456_U.if_full_n;
    assign fifo_intf_1809.fifo_rd_block = 0;
    assign fifo_intf_1809.fifo_wr_block = 0;
    assign fifo_intf_1809.finish = finish;
    csv_file_dump fifo_csv_dumper_1809;
    csv_file_dump cstatus_csv_dumper_1809;
    df_fifo_monitor fifo_monitor_1809;
    df_fifo_intf fifo_intf_1810(clock,reset);
    assign fifo_intf_1810.rd_en = AESL_inst_myproject.layer3_out_457_U.if_read & AESL_inst_myproject.layer3_out_457_U.if_empty_n;
    assign fifo_intf_1810.wr_en = AESL_inst_myproject.layer3_out_457_U.if_write & AESL_inst_myproject.layer3_out_457_U.if_full_n;
    assign fifo_intf_1810.fifo_rd_block = 0;
    assign fifo_intf_1810.fifo_wr_block = 0;
    assign fifo_intf_1810.finish = finish;
    csv_file_dump fifo_csv_dumper_1810;
    csv_file_dump cstatus_csv_dumper_1810;
    df_fifo_monitor fifo_monitor_1810;
    df_fifo_intf fifo_intf_1811(clock,reset);
    assign fifo_intf_1811.rd_en = AESL_inst_myproject.layer3_out_458_U.if_read & AESL_inst_myproject.layer3_out_458_U.if_empty_n;
    assign fifo_intf_1811.wr_en = AESL_inst_myproject.layer3_out_458_U.if_write & AESL_inst_myproject.layer3_out_458_U.if_full_n;
    assign fifo_intf_1811.fifo_rd_block = 0;
    assign fifo_intf_1811.fifo_wr_block = 0;
    assign fifo_intf_1811.finish = finish;
    csv_file_dump fifo_csv_dumper_1811;
    csv_file_dump cstatus_csv_dumper_1811;
    df_fifo_monitor fifo_monitor_1811;
    df_fifo_intf fifo_intf_1812(clock,reset);
    assign fifo_intf_1812.rd_en = AESL_inst_myproject.layer3_out_459_U.if_read & AESL_inst_myproject.layer3_out_459_U.if_empty_n;
    assign fifo_intf_1812.wr_en = AESL_inst_myproject.layer3_out_459_U.if_write & AESL_inst_myproject.layer3_out_459_U.if_full_n;
    assign fifo_intf_1812.fifo_rd_block = 0;
    assign fifo_intf_1812.fifo_wr_block = 0;
    assign fifo_intf_1812.finish = finish;
    csv_file_dump fifo_csv_dumper_1812;
    csv_file_dump cstatus_csv_dumper_1812;
    df_fifo_monitor fifo_monitor_1812;
    df_fifo_intf fifo_intf_1813(clock,reset);
    assign fifo_intf_1813.rd_en = AESL_inst_myproject.layer3_out_460_U.if_read & AESL_inst_myproject.layer3_out_460_U.if_empty_n;
    assign fifo_intf_1813.wr_en = AESL_inst_myproject.layer3_out_460_U.if_write & AESL_inst_myproject.layer3_out_460_U.if_full_n;
    assign fifo_intf_1813.fifo_rd_block = 0;
    assign fifo_intf_1813.fifo_wr_block = 0;
    assign fifo_intf_1813.finish = finish;
    csv_file_dump fifo_csv_dumper_1813;
    csv_file_dump cstatus_csv_dumper_1813;
    df_fifo_monitor fifo_monitor_1813;
    df_fifo_intf fifo_intf_1814(clock,reset);
    assign fifo_intf_1814.rd_en = AESL_inst_myproject.layer3_out_461_U.if_read & AESL_inst_myproject.layer3_out_461_U.if_empty_n;
    assign fifo_intf_1814.wr_en = AESL_inst_myproject.layer3_out_461_U.if_write & AESL_inst_myproject.layer3_out_461_U.if_full_n;
    assign fifo_intf_1814.fifo_rd_block = 0;
    assign fifo_intf_1814.fifo_wr_block = 0;
    assign fifo_intf_1814.finish = finish;
    csv_file_dump fifo_csv_dumper_1814;
    csv_file_dump cstatus_csv_dumper_1814;
    df_fifo_monitor fifo_monitor_1814;
    df_fifo_intf fifo_intf_1815(clock,reset);
    assign fifo_intf_1815.rd_en = AESL_inst_myproject.layer3_out_462_U.if_read & AESL_inst_myproject.layer3_out_462_U.if_empty_n;
    assign fifo_intf_1815.wr_en = AESL_inst_myproject.layer3_out_462_U.if_write & AESL_inst_myproject.layer3_out_462_U.if_full_n;
    assign fifo_intf_1815.fifo_rd_block = 0;
    assign fifo_intf_1815.fifo_wr_block = 0;
    assign fifo_intf_1815.finish = finish;
    csv_file_dump fifo_csv_dumper_1815;
    csv_file_dump cstatus_csv_dumper_1815;
    df_fifo_monitor fifo_monitor_1815;
    df_fifo_intf fifo_intf_1816(clock,reset);
    assign fifo_intf_1816.rd_en = AESL_inst_myproject.layer3_out_463_U.if_read & AESL_inst_myproject.layer3_out_463_U.if_empty_n;
    assign fifo_intf_1816.wr_en = AESL_inst_myproject.layer3_out_463_U.if_write & AESL_inst_myproject.layer3_out_463_U.if_full_n;
    assign fifo_intf_1816.fifo_rd_block = 0;
    assign fifo_intf_1816.fifo_wr_block = 0;
    assign fifo_intf_1816.finish = finish;
    csv_file_dump fifo_csv_dumper_1816;
    csv_file_dump cstatus_csv_dumper_1816;
    df_fifo_monitor fifo_monitor_1816;
    df_fifo_intf fifo_intf_1817(clock,reset);
    assign fifo_intf_1817.rd_en = AESL_inst_myproject.layer3_out_464_U.if_read & AESL_inst_myproject.layer3_out_464_U.if_empty_n;
    assign fifo_intf_1817.wr_en = AESL_inst_myproject.layer3_out_464_U.if_write & AESL_inst_myproject.layer3_out_464_U.if_full_n;
    assign fifo_intf_1817.fifo_rd_block = 0;
    assign fifo_intf_1817.fifo_wr_block = 0;
    assign fifo_intf_1817.finish = finish;
    csv_file_dump fifo_csv_dumper_1817;
    csv_file_dump cstatus_csv_dumper_1817;
    df_fifo_monitor fifo_monitor_1817;
    df_fifo_intf fifo_intf_1818(clock,reset);
    assign fifo_intf_1818.rd_en = AESL_inst_myproject.layer3_out_465_U.if_read & AESL_inst_myproject.layer3_out_465_U.if_empty_n;
    assign fifo_intf_1818.wr_en = AESL_inst_myproject.layer3_out_465_U.if_write & AESL_inst_myproject.layer3_out_465_U.if_full_n;
    assign fifo_intf_1818.fifo_rd_block = 0;
    assign fifo_intf_1818.fifo_wr_block = 0;
    assign fifo_intf_1818.finish = finish;
    csv_file_dump fifo_csv_dumper_1818;
    csv_file_dump cstatus_csv_dumper_1818;
    df_fifo_monitor fifo_monitor_1818;
    df_fifo_intf fifo_intf_1819(clock,reset);
    assign fifo_intf_1819.rd_en = AESL_inst_myproject.layer3_out_466_U.if_read & AESL_inst_myproject.layer3_out_466_U.if_empty_n;
    assign fifo_intf_1819.wr_en = AESL_inst_myproject.layer3_out_466_U.if_write & AESL_inst_myproject.layer3_out_466_U.if_full_n;
    assign fifo_intf_1819.fifo_rd_block = 0;
    assign fifo_intf_1819.fifo_wr_block = 0;
    assign fifo_intf_1819.finish = finish;
    csv_file_dump fifo_csv_dumper_1819;
    csv_file_dump cstatus_csv_dumper_1819;
    df_fifo_monitor fifo_monitor_1819;
    df_fifo_intf fifo_intf_1820(clock,reset);
    assign fifo_intf_1820.rd_en = AESL_inst_myproject.layer3_out_467_U.if_read & AESL_inst_myproject.layer3_out_467_U.if_empty_n;
    assign fifo_intf_1820.wr_en = AESL_inst_myproject.layer3_out_467_U.if_write & AESL_inst_myproject.layer3_out_467_U.if_full_n;
    assign fifo_intf_1820.fifo_rd_block = 0;
    assign fifo_intf_1820.fifo_wr_block = 0;
    assign fifo_intf_1820.finish = finish;
    csv_file_dump fifo_csv_dumper_1820;
    csv_file_dump cstatus_csv_dumper_1820;
    df_fifo_monitor fifo_monitor_1820;
    df_fifo_intf fifo_intf_1821(clock,reset);
    assign fifo_intf_1821.rd_en = AESL_inst_myproject.layer3_out_468_U.if_read & AESL_inst_myproject.layer3_out_468_U.if_empty_n;
    assign fifo_intf_1821.wr_en = AESL_inst_myproject.layer3_out_468_U.if_write & AESL_inst_myproject.layer3_out_468_U.if_full_n;
    assign fifo_intf_1821.fifo_rd_block = 0;
    assign fifo_intf_1821.fifo_wr_block = 0;
    assign fifo_intf_1821.finish = finish;
    csv_file_dump fifo_csv_dumper_1821;
    csv_file_dump cstatus_csv_dumper_1821;
    df_fifo_monitor fifo_monitor_1821;
    df_fifo_intf fifo_intf_1822(clock,reset);
    assign fifo_intf_1822.rd_en = AESL_inst_myproject.layer3_out_469_U.if_read & AESL_inst_myproject.layer3_out_469_U.if_empty_n;
    assign fifo_intf_1822.wr_en = AESL_inst_myproject.layer3_out_469_U.if_write & AESL_inst_myproject.layer3_out_469_U.if_full_n;
    assign fifo_intf_1822.fifo_rd_block = 0;
    assign fifo_intf_1822.fifo_wr_block = 0;
    assign fifo_intf_1822.finish = finish;
    csv_file_dump fifo_csv_dumper_1822;
    csv_file_dump cstatus_csv_dumper_1822;
    df_fifo_monitor fifo_monitor_1822;
    df_fifo_intf fifo_intf_1823(clock,reset);
    assign fifo_intf_1823.rd_en = AESL_inst_myproject.layer3_out_470_U.if_read & AESL_inst_myproject.layer3_out_470_U.if_empty_n;
    assign fifo_intf_1823.wr_en = AESL_inst_myproject.layer3_out_470_U.if_write & AESL_inst_myproject.layer3_out_470_U.if_full_n;
    assign fifo_intf_1823.fifo_rd_block = 0;
    assign fifo_intf_1823.fifo_wr_block = 0;
    assign fifo_intf_1823.finish = finish;
    csv_file_dump fifo_csv_dumper_1823;
    csv_file_dump cstatus_csv_dumper_1823;
    df_fifo_monitor fifo_monitor_1823;
    df_fifo_intf fifo_intf_1824(clock,reset);
    assign fifo_intf_1824.rd_en = AESL_inst_myproject.layer3_out_471_U.if_read & AESL_inst_myproject.layer3_out_471_U.if_empty_n;
    assign fifo_intf_1824.wr_en = AESL_inst_myproject.layer3_out_471_U.if_write & AESL_inst_myproject.layer3_out_471_U.if_full_n;
    assign fifo_intf_1824.fifo_rd_block = 0;
    assign fifo_intf_1824.fifo_wr_block = 0;
    assign fifo_intf_1824.finish = finish;
    csv_file_dump fifo_csv_dumper_1824;
    csv_file_dump cstatus_csv_dumper_1824;
    df_fifo_monitor fifo_monitor_1824;
    df_fifo_intf fifo_intf_1825(clock,reset);
    assign fifo_intf_1825.rd_en = AESL_inst_myproject.layer3_out_472_U.if_read & AESL_inst_myproject.layer3_out_472_U.if_empty_n;
    assign fifo_intf_1825.wr_en = AESL_inst_myproject.layer3_out_472_U.if_write & AESL_inst_myproject.layer3_out_472_U.if_full_n;
    assign fifo_intf_1825.fifo_rd_block = 0;
    assign fifo_intf_1825.fifo_wr_block = 0;
    assign fifo_intf_1825.finish = finish;
    csv_file_dump fifo_csv_dumper_1825;
    csv_file_dump cstatus_csv_dumper_1825;
    df_fifo_monitor fifo_monitor_1825;
    df_fifo_intf fifo_intf_1826(clock,reset);
    assign fifo_intf_1826.rd_en = AESL_inst_myproject.layer3_out_473_U.if_read & AESL_inst_myproject.layer3_out_473_U.if_empty_n;
    assign fifo_intf_1826.wr_en = AESL_inst_myproject.layer3_out_473_U.if_write & AESL_inst_myproject.layer3_out_473_U.if_full_n;
    assign fifo_intf_1826.fifo_rd_block = 0;
    assign fifo_intf_1826.fifo_wr_block = 0;
    assign fifo_intf_1826.finish = finish;
    csv_file_dump fifo_csv_dumper_1826;
    csv_file_dump cstatus_csv_dumper_1826;
    df_fifo_monitor fifo_monitor_1826;
    df_fifo_intf fifo_intf_1827(clock,reset);
    assign fifo_intf_1827.rd_en = AESL_inst_myproject.layer3_out_474_U.if_read & AESL_inst_myproject.layer3_out_474_U.if_empty_n;
    assign fifo_intf_1827.wr_en = AESL_inst_myproject.layer3_out_474_U.if_write & AESL_inst_myproject.layer3_out_474_U.if_full_n;
    assign fifo_intf_1827.fifo_rd_block = 0;
    assign fifo_intf_1827.fifo_wr_block = 0;
    assign fifo_intf_1827.finish = finish;
    csv_file_dump fifo_csv_dumper_1827;
    csv_file_dump cstatus_csv_dumper_1827;
    df_fifo_monitor fifo_monitor_1827;
    df_fifo_intf fifo_intf_1828(clock,reset);
    assign fifo_intf_1828.rd_en = AESL_inst_myproject.layer3_out_475_U.if_read & AESL_inst_myproject.layer3_out_475_U.if_empty_n;
    assign fifo_intf_1828.wr_en = AESL_inst_myproject.layer3_out_475_U.if_write & AESL_inst_myproject.layer3_out_475_U.if_full_n;
    assign fifo_intf_1828.fifo_rd_block = 0;
    assign fifo_intf_1828.fifo_wr_block = 0;
    assign fifo_intf_1828.finish = finish;
    csv_file_dump fifo_csv_dumper_1828;
    csv_file_dump cstatus_csv_dumper_1828;
    df_fifo_monitor fifo_monitor_1828;
    df_fifo_intf fifo_intf_1829(clock,reset);
    assign fifo_intf_1829.rd_en = AESL_inst_myproject.layer3_out_476_U.if_read & AESL_inst_myproject.layer3_out_476_U.if_empty_n;
    assign fifo_intf_1829.wr_en = AESL_inst_myproject.layer3_out_476_U.if_write & AESL_inst_myproject.layer3_out_476_U.if_full_n;
    assign fifo_intf_1829.fifo_rd_block = 0;
    assign fifo_intf_1829.fifo_wr_block = 0;
    assign fifo_intf_1829.finish = finish;
    csv_file_dump fifo_csv_dumper_1829;
    csv_file_dump cstatus_csv_dumper_1829;
    df_fifo_monitor fifo_monitor_1829;
    df_fifo_intf fifo_intf_1830(clock,reset);
    assign fifo_intf_1830.rd_en = AESL_inst_myproject.layer3_out_477_U.if_read & AESL_inst_myproject.layer3_out_477_U.if_empty_n;
    assign fifo_intf_1830.wr_en = AESL_inst_myproject.layer3_out_477_U.if_write & AESL_inst_myproject.layer3_out_477_U.if_full_n;
    assign fifo_intf_1830.fifo_rd_block = 0;
    assign fifo_intf_1830.fifo_wr_block = 0;
    assign fifo_intf_1830.finish = finish;
    csv_file_dump fifo_csv_dumper_1830;
    csv_file_dump cstatus_csv_dumper_1830;
    df_fifo_monitor fifo_monitor_1830;
    df_fifo_intf fifo_intf_1831(clock,reset);
    assign fifo_intf_1831.rd_en = AESL_inst_myproject.layer3_out_478_U.if_read & AESL_inst_myproject.layer3_out_478_U.if_empty_n;
    assign fifo_intf_1831.wr_en = AESL_inst_myproject.layer3_out_478_U.if_write & AESL_inst_myproject.layer3_out_478_U.if_full_n;
    assign fifo_intf_1831.fifo_rd_block = 0;
    assign fifo_intf_1831.fifo_wr_block = 0;
    assign fifo_intf_1831.finish = finish;
    csv_file_dump fifo_csv_dumper_1831;
    csv_file_dump cstatus_csv_dumper_1831;
    df_fifo_monitor fifo_monitor_1831;
    df_fifo_intf fifo_intf_1832(clock,reset);
    assign fifo_intf_1832.rd_en = AESL_inst_myproject.layer3_out_479_U.if_read & AESL_inst_myproject.layer3_out_479_U.if_empty_n;
    assign fifo_intf_1832.wr_en = AESL_inst_myproject.layer3_out_479_U.if_write & AESL_inst_myproject.layer3_out_479_U.if_full_n;
    assign fifo_intf_1832.fifo_rd_block = 0;
    assign fifo_intf_1832.fifo_wr_block = 0;
    assign fifo_intf_1832.finish = finish;
    csv_file_dump fifo_csv_dumper_1832;
    csv_file_dump cstatus_csv_dumper_1832;
    df_fifo_monitor fifo_monitor_1832;
    df_fifo_intf fifo_intf_1833(clock,reset);
    assign fifo_intf_1833.rd_en = AESL_inst_myproject.layer3_out_480_U.if_read & AESL_inst_myproject.layer3_out_480_U.if_empty_n;
    assign fifo_intf_1833.wr_en = AESL_inst_myproject.layer3_out_480_U.if_write & AESL_inst_myproject.layer3_out_480_U.if_full_n;
    assign fifo_intf_1833.fifo_rd_block = 0;
    assign fifo_intf_1833.fifo_wr_block = 0;
    assign fifo_intf_1833.finish = finish;
    csv_file_dump fifo_csv_dumper_1833;
    csv_file_dump cstatus_csv_dumper_1833;
    df_fifo_monitor fifo_monitor_1833;
    df_fifo_intf fifo_intf_1834(clock,reset);
    assign fifo_intf_1834.rd_en = AESL_inst_myproject.layer3_out_481_U.if_read & AESL_inst_myproject.layer3_out_481_U.if_empty_n;
    assign fifo_intf_1834.wr_en = AESL_inst_myproject.layer3_out_481_U.if_write & AESL_inst_myproject.layer3_out_481_U.if_full_n;
    assign fifo_intf_1834.fifo_rd_block = 0;
    assign fifo_intf_1834.fifo_wr_block = 0;
    assign fifo_intf_1834.finish = finish;
    csv_file_dump fifo_csv_dumper_1834;
    csv_file_dump cstatus_csv_dumper_1834;
    df_fifo_monitor fifo_monitor_1834;
    df_fifo_intf fifo_intf_1835(clock,reset);
    assign fifo_intf_1835.rd_en = AESL_inst_myproject.layer3_out_482_U.if_read & AESL_inst_myproject.layer3_out_482_U.if_empty_n;
    assign fifo_intf_1835.wr_en = AESL_inst_myproject.layer3_out_482_U.if_write & AESL_inst_myproject.layer3_out_482_U.if_full_n;
    assign fifo_intf_1835.fifo_rd_block = 0;
    assign fifo_intf_1835.fifo_wr_block = 0;
    assign fifo_intf_1835.finish = finish;
    csv_file_dump fifo_csv_dumper_1835;
    csv_file_dump cstatus_csv_dumper_1835;
    df_fifo_monitor fifo_monitor_1835;
    df_fifo_intf fifo_intf_1836(clock,reset);
    assign fifo_intf_1836.rd_en = AESL_inst_myproject.layer3_out_483_U.if_read & AESL_inst_myproject.layer3_out_483_U.if_empty_n;
    assign fifo_intf_1836.wr_en = AESL_inst_myproject.layer3_out_483_U.if_write & AESL_inst_myproject.layer3_out_483_U.if_full_n;
    assign fifo_intf_1836.fifo_rd_block = 0;
    assign fifo_intf_1836.fifo_wr_block = 0;
    assign fifo_intf_1836.finish = finish;
    csv_file_dump fifo_csv_dumper_1836;
    csv_file_dump cstatus_csv_dumper_1836;
    df_fifo_monitor fifo_monitor_1836;
    df_fifo_intf fifo_intf_1837(clock,reset);
    assign fifo_intf_1837.rd_en = AESL_inst_myproject.layer3_out_484_U.if_read & AESL_inst_myproject.layer3_out_484_U.if_empty_n;
    assign fifo_intf_1837.wr_en = AESL_inst_myproject.layer3_out_484_U.if_write & AESL_inst_myproject.layer3_out_484_U.if_full_n;
    assign fifo_intf_1837.fifo_rd_block = 0;
    assign fifo_intf_1837.fifo_wr_block = 0;
    assign fifo_intf_1837.finish = finish;
    csv_file_dump fifo_csv_dumper_1837;
    csv_file_dump cstatus_csv_dumper_1837;
    df_fifo_monitor fifo_monitor_1837;
    df_fifo_intf fifo_intf_1838(clock,reset);
    assign fifo_intf_1838.rd_en = AESL_inst_myproject.layer3_out_485_U.if_read & AESL_inst_myproject.layer3_out_485_U.if_empty_n;
    assign fifo_intf_1838.wr_en = AESL_inst_myproject.layer3_out_485_U.if_write & AESL_inst_myproject.layer3_out_485_U.if_full_n;
    assign fifo_intf_1838.fifo_rd_block = 0;
    assign fifo_intf_1838.fifo_wr_block = 0;
    assign fifo_intf_1838.finish = finish;
    csv_file_dump fifo_csv_dumper_1838;
    csv_file_dump cstatus_csv_dumper_1838;
    df_fifo_monitor fifo_monitor_1838;
    df_fifo_intf fifo_intf_1839(clock,reset);
    assign fifo_intf_1839.rd_en = AESL_inst_myproject.layer3_out_486_U.if_read & AESL_inst_myproject.layer3_out_486_U.if_empty_n;
    assign fifo_intf_1839.wr_en = AESL_inst_myproject.layer3_out_486_U.if_write & AESL_inst_myproject.layer3_out_486_U.if_full_n;
    assign fifo_intf_1839.fifo_rd_block = 0;
    assign fifo_intf_1839.fifo_wr_block = 0;
    assign fifo_intf_1839.finish = finish;
    csv_file_dump fifo_csv_dumper_1839;
    csv_file_dump cstatus_csv_dumper_1839;
    df_fifo_monitor fifo_monitor_1839;
    df_fifo_intf fifo_intf_1840(clock,reset);
    assign fifo_intf_1840.rd_en = AESL_inst_myproject.layer3_out_487_U.if_read & AESL_inst_myproject.layer3_out_487_U.if_empty_n;
    assign fifo_intf_1840.wr_en = AESL_inst_myproject.layer3_out_487_U.if_write & AESL_inst_myproject.layer3_out_487_U.if_full_n;
    assign fifo_intf_1840.fifo_rd_block = 0;
    assign fifo_intf_1840.fifo_wr_block = 0;
    assign fifo_intf_1840.finish = finish;
    csv_file_dump fifo_csv_dumper_1840;
    csv_file_dump cstatus_csv_dumper_1840;
    df_fifo_monitor fifo_monitor_1840;
    df_fifo_intf fifo_intf_1841(clock,reset);
    assign fifo_intf_1841.rd_en = AESL_inst_myproject.layer3_out_488_U.if_read & AESL_inst_myproject.layer3_out_488_U.if_empty_n;
    assign fifo_intf_1841.wr_en = AESL_inst_myproject.layer3_out_488_U.if_write & AESL_inst_myproject.layer3_out_488_U.if_full_n;
    assign fifo_intf_1841.fifo_rd_block = 0;
    assign fifo_intf_1841.fifo_wr_block = 0;
    assign fifo_intf_1841.finish = finish;
    csv_file_dump fifo_csv_dumper_1841;
    csv_file_dump cstatus_csv_dumper_1841;
    df_fifo_monitor fifo_monitor_1841;
    df_fifo_intf fifo_intf_1842(clock,reset);
    assign fifo_intf_1842.rd_en = AESL_inst_myproject.layer3_out_489_U.if_read & AESL_inst_myproject.layer3_out_489_U.if_empty_n;
    assign fifo_intf_1842.wr_en = AESL_inst_myproject.layer3_out_489_U.if_write & AESL_inst_myproject.layer3_out_489_U.if_full_n;
    assign fifo_intf_1842.fifo_rd_block = 0;
    assign fifo_intf_1842.fifo_wr_block = 0;
    assign fifo_intf_1842.finish = finish;
    csv_file_dump fifo_csv_dumper_1842;
    csv_file_dump cstatus_csv_dumper_1842;
    df_fifo_monitor fifo_monitor_1842;
    df_fifo_intf fifo_intf_1843(clock,reset);
    assign fifo_intf_1843.rd_en = AESL_inst_myproject.layer3_out_490_U.if_read & AESL_inst_myproject.layer3_out_490_U.if_empty_n;
    assign fifo_intf_1843.wr_en = AESL_inst_myproject.layer3_out_490_U.if_write & AESL_inst_myproject.layer3_out_490_U.if_full_n;
    assign fifo_intf_1843.fifo_rd_block = 0;
    assign fifo_intf_1843.fifo_wr_block = 0;
    assign fifo_intf_1843.finish = finish;
    csv_file_dump fifo_csv_dumper_1843;
    csv_file_dump cstatus_csv_dumper_1843;
    df_fifo_monitor fifo_monitor_1843;
    df_fifo_intf fifo_intf_1844(clock,reset);
    assign fifo_intf_1844.rd_en = AESL_inst_myproject.layer3_out_491_U.if_read & AESL_inst_myproject.layer3_out_491_U.if_empty_n;
    assign fifo_intf_1844.wr_en = AESL_inst_myproject.layer3_out_491_U.if_write & AESL_inst_myproject.layer3_out_491_U.if_full_n;
    assign fifo_intf_1844.fifo_rd_block = 0;
    assign fifo_intf_1844.fifo_wr_block = 0;
    assign fifo_intf_1844.finish = finish;
    csv_file_dump fifo_csv_dumper_1844;
    csv_file_dump cstatus_csv_dumper_1844;
    df_fifo_monitor fifo_monitor_1844;
    df_fifo_intf fifo_intf_1845(clock,reset);
    assign fifo_intf_1845.rd_en = AESL_inst_myproject.layer3_out_492_U.if_read & AESL_inst_myproject.layer3_out_492_U.if_empty_n;
    assign fifo_intf_1845.wr_en = AESL_inst_myproject.layer3_out_492_U.if_write & AESL_inst_myproject.layer3_out_492_U.if_full_n;
    assign fifo_intf_1845.fifo_rd_block = 0;
    assign fifo_intf_1845.fifo_wr_block = 0;
    assign fifo_intf_1845.finish = finish;
    csv_file_dump fifo_csv_dumper_1845;
    csv_file_dump cstatus_csv_dumper_1845;
    df_fifo_monitor fifo_monitor_1845;
    df_fifo_intf fifo_intf_1846(clock,reset);
    assign fifo_intf_1846.rd_en = AESL_inst_myproject.layer3_out_493_U.if_read & AESL_inst_myproject.layer3_out_493_U.if_empty_n;
    assign fifo_intf_1846.wr_en = AESL_inst_myproject.layer3_out_493_U.if_write & AESL_inst_myproject.layer3_out_493_U.if_full_n;
    assign fifo_intf_1846.fifo_rd_block = 0;
    assign fifo_intf_1846.fifo_wr_block = 0;
    assign fifo_intf_1846.finish = finish;
    csv_file_dump fifo_csv_dumper_1846;
    csv_file_dump cstatus_csv_dumper_1846;
    df_fifo_monitor fifo_monitor_1846;
    df_fifo_intf fifo_intf_1847(clock,reset);
    assign fifo_intf_1847.rd_en = AESL_inst_myproject.layer3_out_494_U.if_read & AESL_inst_myproject.layer3_out_494_U.if_empty_n;
    assign fifo_intf_1847.wr_en = AESL_inst_myproject.layer3_out_494_U.if_write & AESL_inst_myproject.layer3_out_494_U.if_full_n;
    assign fifo_intf_1847.fifo_rd_block = 0;
    assign fifo_intf_1847.fifo_wr_block = 0;
    assign fifo_intf_1847.finish = finish;
    csv_file_dump fifo_csv_dumper_1847;
    csv_file_dump cstatus_csv_dumper_1847;
    df_fifo_monitor fifo_monitor_1847;
    df_fifo_intf fifo_intf_1848(clock,reset);
    assign fifo_intf_1848.rd_en = AESL_inst_myproject.layer3_out_495_U.if_read & AESL_inst_myproject.layer3_out_495_U.if_empty_n;
    assign fifo_intf_1848.wr_en = AESL_inst_myproject.layer3_out_495_U.if_write & AESL_inst_myproject.layer3_out_495_U.if_full_n;
    assign fifo_intf_1848.fifo_rd_block = 0;
    assign fifo_intf_1848.fifo_wr_block = 0;
    assign fifo_intf_1848.finish = finish;
    csv_file_dump fifo_csv_dumper_1848;
    csv_file_dump cstatus_csv_dumper_1848;
    df_fifo_monitor fifo_monitor_1848;
    df_fifo_intf fifo_intf_1849(clock,reset);
    assign fifo_intf_1849.rd_en = AESL_inst_myproject.layer3_out_496_U.if_read & AESL_inst_myproject.layer3_out_496_U.if_empty_n;
    assign fifo_intf_1849.wr_en = AESL_inst_myproject.layer3_out_496_U.if_write & AESL_inst_myproject.layer3_out_496_U.if_full_n;
    assign fifo_intf_1849.fifo_rd_block = 0;
    assign fifo_intf_1849.fifo_wr_block = 0;
    assign fifo_intf_1849.finish = finish;
    csv_file_dump fifo_csv_dumper_1849;
    csv_file_dump cstatus_csv_dumper_1849;
    df_fifo_monitor fifo_monitor_1849;
    df_fifo_intf fifo_intf_1850(clock,reset);
    assign fifo_intf_1850.rd_en = AESL_inst_myproject.layer3_out_497_U.if_read & AESL_inst_myproject.layer3_out_497_U.if_empty_n;
    assign fifo_intf_1850.wr_en = AESL_inst_myproject.layer3_out_497_U.if_write & AESL_inst_myproject.layer3_out_497_U.if_full_n;
    assign fifo_intf_1850.fifo_rd_block = 0;
    assign fifo_intf_1850.fifo_wr_block = 0;
    assign fifo_intf_1850.finish = finish;
    csv_file_dump fifo_csv_dumper_1850;
    csv_file_dump cstatus_csv_dumper_1850;
    df_fifo_monitor fifo_monitor_1850;
    df_fifo_intf fifo_intf_1851(clock,reset);
    assign fifo_intf_1851.rd_en = AESL_inst_myproject.layer3_out_498_U.if_read & AESL_inst_myproject.layer3_out_498_U.if_empty_n;
    assign fifo_intf_1851.wr_en = AESL_inst_myproject.layer3_out_498_U.if_write & AESL_inst_myproject.layer3_out_498_U.if_full_n;
    assign fifo_intf_1851.fifo_rd_block = 0;
    assign fifo_intf_1851.fifo_wr_block = 0;
    assign fifo_intf_1851.finish = finish;
    csv_file_dump fifo_csv_dumper_1851;
    csv_file_dump cstatus_csv_dumper_1851;
    df_fifo_monitor fifo_monitor_1851;
    df_fifo_intf fifo_intf_1852(clock,reset);
    assign fifo_intf_1852.rd_en = AESL_inst_myproject.layer3_out_499_U.if_read & AESL_inst_myproject.layer3_out_499_U.if_empty_n;
    assign fifo_intf_1852.wr_en = AESL_inst_myproject.layer3_out_499_U.if_write & AESL_inst_myproject.layer3_out_499_U.if_full_n;
    assign fifo_intf_1852.fifo_rd_block = 0;
    assign fifo_intf_1852.fifo_wr_block = 0;
    assign fifo_intf_1852.finish = finish;
    csv_file_dump fifo_csv_dumper_1852;
    csv_file_dump cstatus_csv_dumper_1852;
    df_fifo_monitor fifo_monitor_1852;
    df_fifo_intf fifo_intf_1853(clock,reset);
    assign fifo_intf_1853.rd_en = AESL_inst_myproject.layer3_out_500_U.if_read & AESL_inst_myproject.layer3_out_500_U.if_empty_n;
    assign fifo_intf_1853.wr_en = AESL_inst_myproject.layer3_out_500_U.if_write & AESL_inst_myproject.layer3_out_500_U.if_full_n;
    assign fifo_intf_1853.fifo_rd_block = 0;
    assign fifo_intf_1853.fifo_wr_block = 0;
    assign fifo_intf_1853.finish = finish;
    csv_file_dump fifo_csv_dumper_1853;
    csv_file_dump cstatus_csv_dumper_1853;
    df_fifo_monitor fifo_monitor_1853;
    df_fifo_intf fifo_intf_1854(clock,reset);
    assign fifo_intf_1854.rd_en = AESL_inst_myproject.layer3_out_501_U.if_read & AESL_inst_myproject.layer3_out_501_U.if_empty_n;
    assign fifo_intf_1854.wr_en = AESL_inst_myproject.layer3_out_501_U.if_write & AESL_inst_myproject.layer3_out_501_U.if_full_n;
    assign fifo_intf_1854.fifo_rd_block = 0;
    assign fifo_intf_1854.fifo_wr_block = 0;
    assign fifo_intf_1854.finish = finish;
    csv_file_dump fifo_csv_dumper_1854;
    csv_file_dump cstatus_csv_dumper_1854;
    df_fifo_monitor fifo_monitor_1854;
    df_fifo_intf fifo_intf_1855(clock,reset);
    assign fifo_intf_1855.rd_en = AESL_inst_myproject.layer3_out_502_U.if_read & AESL_inst_myproject.layer3_out_502_U.if_empty_n;
    assign fifo_intf_1855.wr_en = AESL_inst_myproject.layer3_out_502_U.if_write & AESL_inst_myproject.layer3_out_502_U.if_full_n;
    assign fifo_intf_1855.fifo_rd_block = 0;
    assign fifo_intf_1855.fifo_wr_block = 0;
    assign fifo_intf_1855.finish = finish;
    csv_file_dump fifo_csv_dumper_1855;
    csv_file_dump cstatus_csv_dumper_1855;
    df_fifo_monitor fifo_monitor_1855;
    df_fifo_intf fifo_intf_1856(clock,reset);
    assign fifo_intf_1856.rd_en = AESL_inst_myproject.layer3_out_503_U.if_read & AESL_inst_myproject.layer3_out_503_U.if_empty_n;
    assign fifo_intf_1856.wr_en = AESL_inst_myproject.layer3_out_503_U.if_write & AESL_inst_myproject.layer3_out_503_U.if_full_n;
    assign fifo_intf_1856.fifo_rd_block = 0;
    assign fifo_intf_1856.fifo_wr_block = 0;
    assign fifo_intf_1856.finish = finish;
    csv_file_dump fifo_csv_dumper_1856;
    csv_file_dump cstatus_csv_dumper_1856;
    df_fifo_monitor fifo_monitor_1856;
    df_fifo_intf fifo_intf_1857(clock,reset);
    assign fifo_intf_1857.rd_en = AESL_inst_myproject.layer3_out_504_U.if_read & AESL_inst_myproject.layer3_out_504_U.if_empty_n;
    assign fifo_intf_1857.wr_en = AESL_inst_myproject.layer3_out_504_U.if_write & AESL_inst_myproject.layer3_out_504_U.if_full_n;
    assign fifo_intf_1857.fifo_rd_block = 0;
    assign fifo_intf_1857.fifo_wr_block = 0;
    assign fifo_intf_1857.finish = finish;
    csv_file_dump fifo_csv_dumper_1857;
    csv_file_dump cstatus_csv_dumper_1857;
    df_fifo_monitor fifo_monitor_1857;
    df_fifo_intf fifo_intf_1858(clock,reset);
    assign fifo_intf_1858.rd_en = AESL_inst_myproject.layer3_out_505_U.if_read & AESL_inst_myproject.layer3_out_505_U.if_empty_n;
    assign fifo_intf_1858.wr_en = AESL_inst_myproject.layer3_out_505_U.if_write & AESL_inst_myproject.layer3_out_505_U.if_full_n;
    assign fifo_intf_1858.fifo_rd_block = 0;
    assign fifo_intf_1858.fifo_wr_block = 0;
    assign fifo_intf_1858.finish = finish;
    csv_file_dump fifo_csv_dumper_1858;
    csv_file_dump cstatus_csv_dumper_1858;
    df_fifo_monitor fifo_monitor_1858;
    df_fifo_intf fifo_intf_1859(clock,reset);
    assign fifo_intf_1859.rd_en = AESL_inst_myproject.layer3_out_506_U.if_read & AESL_inst_myproject.layer3_out_506_U.if_empty_n;
    assign fifo_intf_1859.wr_en = AESL_inst_myproject.layer3_out_506_U.if_write & AESL_inst_myproject.layer3_out_506_U.if_full_n;
    assign fifo_intf_1859.fifo_rd_block = 0;
    assign fifo_intf_1859.fifo_wr_block = 0;
    assign fifo_intf_1859.finish = finish;
    csv_file_dump fifo_csv_dumper_1859;
    csv_file_dump cstatus_csv_dumper_1859;
    df_fifo_monitor fifo_monitor_1859;
    df_fifo_intf fifo_intf_1860(clock,reset);
    assign fifo_intf_1860.rd_en = AESL_inst_myproject.layer3_out_507_U.if_read & AESL_inst_myproject.layer3_out_507_U.if_empty_n;
    assign fifo_intf_1860.wr_en = AESL_inst_myproject.layer3_out_507_U.if_write & AESL_inst_myproject.layer3_out_507_U.if_full_n;
    assign fifo_intf_1860.fifo_rd_block = 0;
    assign fifo_intf_1860.fifo_wr_block = 0;
    assign fifo_intf_1860.finish = finish;
    csv_file_dump fifo_csv_dumper_1860;
    csv_file_dump cstatus_csv_dumper_1860;
    df_fifo_monitor fifo_monitor_1860;
    df_fifo_intf fifo_intf_1861(clock,reset);
    assign fifo_intf_1861.rd_en = AESL_inst_myproject.layer3_out_508_U.if_read & AESL_inst_myproject.layer3_out_508_U.if_empty_n;
    assign fifo_intf_1861.wr_en = AESL_inst_myproject.layer3_out_508_U.if_write & AESL_inst_myproject.layer3_out_508_U.if_full_n;
    assign fifo_intf_1861.fifo_rd_block = 0;
    assign fifo_intf_1861.fifo_wr_block = 0;
    assign fifo_intf_1861.finish = finish;
    csv_file_dump fifo_csv_dumper_1861;
    csv_file_dump cstatus_csv_dumper_1861;
    df_fifo_monitor fifo_monitor_1861;
    df_fifo_intf fifo_intf_1862(clock,reset);
    assign fifo_intf_1862.rd_en = AESL_inst_myproject.layer3_out_509_U.if_read & AESL_inst_myproject.layer3_out_509_U.if_empty_n;
    assign fifo_intf_1862.wr_en = AESL_inst_myproject.layer3_out_509_U.if_write & AESL_inst_myproject.layer3_out_509_U.if_full_n;
    assign fifo_intf_1862.fifo_rd_block = 0;
    assign fifo_intf_1862.fifo_wr_block = 0;
    assign fifo_intf_1862.finish = finish;
    csv_file_dump fifo_csv_dumper_1862;
    csv_file_dump cstatus_csv_dumper_1862;
    df_fifo_monitor fifo_monitor_1862;
    df_fifo_intf fifo_intf_1863(clock,reset);
    assign fifo_intf_1863.rd_en = AESL_inst_myproject.layer3_out_510_U.if_read & AESL_inst_myproject.layer3_out_510_U.if_empty_n;
    assign fifo_intf_1863.wr_en = AESL_inst_myproject.layer3_out_510_U.if_write & AESL_inst_myproject.layer3_out_510_U.if_full_n;
    assign fifo_intf_1863.fifo_rd_block = 0;
    assign fifo_intf_1863.fifo_wr_block = 0;
    assign fifo_intf_1863.finish = finish;
    csv_file_dump fifo_csv_dumper_1863;
    csv_file_dump cstatus_csv_dumper_1863;
    df_fifo_monitor fifo_monitor_1863;
    df_fifo_intf fifo_intf_1864(clock,reset);
    assign fifo_intf_1864.rd_en = AESL_inst_myproject.layer3_out_511_U.if_read & AESL_inst_myproject.layer3_out_511_U.if_empty_n;
    assign fifo_intf_1864.wr_en = AESL_inst_myproject.layer3_out_511_U.if_write & AESL_inst_myproject.layer3_out_511_U.if_full_n;
    assign fifo_intf_1864.fifo_rd_block = 0;
    assign fifo_intf_1864.fifo_wr_block = 0;
    assign fifo_intf_1864.finish = finish;
    csv_file_dump fifo_csv_dumper_1864;
    csv_file_dump cstatus_csv_dumper_1864;
    df_fifo_monitor fifo_monitor_1864;
    df_fifo_intf fifo_intf_1865(clock,reset);
    assign fifo_intf_1865.rd_en = AESL_inst_myproject.layer3_out_512_U.if_read & AESL_inst_myproject.layer3_out_512_U.if_empty_n;
    assign fifo_intf_1865.wr_en = AESL_inst_myproject.layer3_out_512_U.if_write & AESL_inst_myproject.layer3_out_512_U.if_full_n;
    assign fifo_intf_1865.fifo_rd_block = 0;
    assign fifo_intf_1865.fifo_wr_block = 0;
    assign fifo_intf_1865.finish = finish;
    csv_file_dump fifo_csv_dumper_1865;
    csv_file_dump cstatus_csv_dumper_1865;
    df_fifo_monitor fifo_monitor_1865;
    df_fifo_intf fifo_intf_1866(clock,reset);
    assign fifo_intf_1866.rd_en = AESL_inst_myproject.layer3_out_513_U.if_read & AESL_inst_myproject.layer3_out_513_U.if_empty_n;
    assign fifo_intf_1866.wr_en = AESL_inst_myproject.layer3_out_513_U.if_write & AESL_inst_myproject.layer3_out_513_U.if_full_n;
    assign fifo_intf_1866.fifo_rd_block = 0;
    assign fifo_intf_1866.fifo_wr_block = 0;
    assign fifo_intf_1866.finish = finish;
    csv_file_dump fifo_csv_dumper_1866;
    csv_file_dump cstatus_csv_dumper_1866;
    df_fifo_monitor fifo_monitor_1866;
    df_fifo_intf fifo_intf_1867(clock,reset);
    assign fifo_intf_1867.rd_en = AESL_inst_myproject.layer3_out_514_U.if_read & AESL_inst_myproject.layer3_out_514_U.if_empty_n;
    assign fifo_intf_1867.wr_en = AESL_inst_myproject.layer3_out_514_U.if_write & AESL_inst_myproject.layer3_out_514_U.if_full_n;
    assign fifo_intf_1867.fifo_rd_block = 0;
    assign fifo_intf_1867.fifo_wr_block = 0;
    assign fifo_intf_1867.finish = finish;
    csv_file_dump fifo_csv_dumper_1867;
    csv_file_dump cstatus_csv_dumper_1867;
    df_fifo_monitor fifo_monitor_1867;
    df_fifo_intf fifo_intf_1868(clock,reset);
    assign fifo_intf_1868.rd_en = AESL_inst_myproject.layer3_out_515_U.if_read & AESL_inst_myproject.layer3_out_515_U.if_empty_n;
    assign fifo_intf_1868.wr_en = AESL_inst_myproject.layer3_out_515_U.if_write & AESL_inst_myproject.layer3_out_515_U.if_full_n;
    assign fifo_intf_1868.fifo_rd_block = 0;
    assign fifo_intf_1868.fifo_wr_block = 0;
    assign fifo_intf_1868.finish = finish;
    csv_file_dump fifo_csv_dumper_1868;
    csv_file_dump cstatus_csv_dumper_1868;
    df_fifo_monitor fifo_monitor_1868;
    df_fifo_intf fifo_intf_1869(clock,reset);
    assign fifo_intf_1869.rd_en = AESL_inst_myproject.layer3_out_516_U.if_read & AESL_inst_myproject.layer3_out_516_U.if_empty_n;
    assign fifo_intf_1869.wr_en = AESL_inst_myproject.layer3_out_516_U.if_write & AESL_inst_myproject.layer3_out_516_U.if_full_n;
    assign fifo_intf_1869.fifo_rd_block = 0;
    assign fifo_intf_1869.fifo_wr_block = 0;
    assign fifo_intf_1869.finish = finish;
    csv_file_dump fifo_csv_dumper_1869;
    csv_file_dump cstatus_csv_dumper_1869;
    df_fifo_monitor fifo_monitor_1869;
    df_fifo_intf fifo_intf_1870(clock,reset);
    assign fifo_intf_1870.rd_en = AESL_inst_myproject.layer3_out_517_U.if_read & AESL_inst_myproject.layer3_out_517_U.if_empty_n;
    assign fifo_intf_1870.wr_en = AESL_inst_myproject.layer3_out_517_U.if_write & AESL_inst_myproject.layer3_out_517_U.if_full_n;
    assign fifo_intf_1870.fifo_rd_block = 0;
    assign fifo_intf_1870.fifo_wr_block = 0;
    assign fifo_intf_1870.finish = finish;
    csv_file_dump fifo_csv_dumper_1870;
    csv_file_dump cstatus_csv_dumper_1870;
    df_fifo_monitor fifo_monitor_1870;
    df_fifo_intf fifo_intf_1871(clock,reset);
    assign fifo_intf_1871.rd_en = AESL_inst_myproject.layer3_out_518_U.if_read & AESL_inst_myproject.layer3_out_518_U.if_empty_n;
    assign fifo_intf_1871.wr_en = AESL_inst_myproject.layer3_out_518_U.if_write & AESL_inst_myproject.layer3_out_518_U.if_full_n;
    assign fifo_intf_1871.fifo_rd_block = 0;
    assign fifo_intf_1871.fifo_wr_block = 0;
    assign fifo_intf_1871.finish = finish;
    csv_file_dump fifo_csv_dumper_1871;
    csv_file_dump cstatus_csv_dumper_1871;
    df_fifo_monitor fifo_monitor_1871;
    df_fifo_intf fifo_intf_1872(clock,reset);
    assign fifo_intf_1872.rd_en = AESL_inst_myproject.layer3_out_519_U.if_read & AESL_inst_myproject.layer3_out_519_U.if_empty_n;
    assign fifo_intf_1872.wr_en = AESL_inst_myproject.layer3_out_519_U.if_write & AESL_inst_myproject.layer3_out_519_U.if_full_n;
    assign fifo_intf_1872.fifo_rd_block = 0;
    assign fifo_intf_1872.fifo_wr_block = 0;
    assign fifo_intf_1872.finish = finish;
    csv_file_dump fifo_csv_dumper_1872;
    csv_file_dump cstatus_csv_dumper_1872;
    df_fifo_monitor fifo_monitor_1872;
    df_fifo_intf fifo_intf_1873(clock,reset);
    assign fifo_intf_1873.rd_en = AESL_inst_myproject.layer3_out_520_U.if_read & AESL_inst_myproject.layer3_out_520_U.if_empty_n;
    assign fifo_intf_1873.wr_en = AESL_inst_myproject.layer3_out_520_U.if_write & AESL_inst_myproject.layer3_out_520_U.if_full_n;
    assign fifo_intf_1873.fifo_rd_block = 0;
    assign fifo_intf_1873.fifo_wr_block = 0;
    assign fifo_intf_1873.finish = finish;
    csv_file_dump fifo_csv_dumper_1873;
    csv_file_dump cstatus_csv_dumper_1873;
    df_fifo_monitor fifo_monitor_1873;
    df_fifo_intf fifo_intf_1874(clock,reset);
    assign fifo_intf_1874.rd_en = AESL_inst_myproject.layer3_out_521_U.if_read & AESL_inst_myproject.layer3_out_521_U.if_empty_n;
    assign fifo_intf_1874.wr_en = AESL_inst_myproject.layer3_out_521_U.if_write & AESL_inst_myproject.layer3_out_521_U.if_full_n;
    assign fifo_intf_1874.fifo_rd_block = 0;
    assign fifo_intf_1874.fifo_wr_block = 0;
    assign fifo_intf_1874.finish = finish;
    csv_file_dump fifo_csv_dumper_1874;
    csv_file_dump cstatus_csv_dumper_1874;
    df_fifo_monitor fifo_monitor_1874;
    df_fifo_intf fifo_intf_1875(clock,reset);
    assign fifo_intf_1875.rd_en = AESL_inst_myproject.layer3_out_522_U.if_read & AESL_inst_myproject.layer3_out_522_U.if_empty_n;
    assign fifo_intf_1875.wr_en = AESL_inst_myproject.layer3_out_522_U.if_write & AESL_inst_myproject.layer3_out_522_U.if_full_n;
    assign fifo_intf_1875.fifo_rd_block = 0;
    assign fifo_intf_1875.fifo_wr_block = 0;
    assign fifo_intf_1875.finish = finish;
    csv_file_dump fifo_csv_dumper_1875;
    csv_file_dump cstatus_csv_dumper_1875;
    df_fifo_monitor fifo_monitor_1875;
    df_fifo_intf fifo_intf_1876(clock,reset);
    assign fifo_intf_1876.rd_en = AESL_inst_myproject.layer3_out_523_U.if_read & AESL_inst_myproject.layer3_out_523_U.if_empty_n;
    assign fifo_intf_1876.wr_en = AESL_inst_myproject.layer3_out_523_U.if_write & AESL_inst_myproject.layer3_out_523_U.if_full_n;
    assign fifo_intf_1876.fifo_rd_block = 0;
    assign fifo_intf_1876.fifo_wr_block = 0;
    assign fifo_intf_1876.finish = finish;
    csv_file_dump fifo_csv_dumper_1876;
    csv_file_dump cstatus_csv_dumper_1876;
    df_fifo_monitor fifo_monitor_1876;
    df_fifo_intf fifo_intf_1877(clock,reset);
    assign fifo_intf_1877.rd_en = AESL_inst_myproject.layer3_out_524_U.if_read & AESL_inst_myproject.layer3_out_524_U.if_empty_n;
    assign fifo_intf_1877.wr_en = AESL_inst_myproject.layer3_out_524_U.if_write & AESL_inst_myproject.layer3_out_524_U.if_full_n;
    assign fifo_intf_1877.fifo_rd_block = 0;
    assign fifo_intf_1877.fifo_wr_block = 0;
    assign fifo_intf_1877.finish = finish;
    csv_file_dump fifo_csv_dumper_1877;
    csv_file_dump cstatus_csv_dumper_1877;
    df_fifo_monitor fifo_monitor_1877;
    df_fifo_intf fifo_intf_1878(clock,reset);
    assign fifo_intf_1878.rd_en = AESL_inst_myproject.layer3_out_525_U.if_read & AESL_inst_myproject.layer3_out_525_U.if_empty_n;
    assign fifo_intf_1878.wr_en = AESL_inst_myproject.layer3_out_525_U.if_write & AESL_inst_myproject.layer3_out_525_U.if_full_n;
    assign fifo_intf_1878.fifo_rd_block = 0;
    assign fifo_intf_1878.fifo_wr_block = 0;
    assign fifo_intf_1878.finish = finish;
    csv_file_dump fifo_csv_dumper_1878;
    csv_file_dump cstatus_csv_dumper_1878;
    df_fifo_monitor fifo_monitor_1878;
    df_fifo_intf fifo_intf_1879(clock,reset);
    assign fifo_intf_1879.rd_en = AESL_inst_myproject.layer3_out_526_U.if_read & AESL_inst_myproject.layer3_out_526_U.if_empty_n;
    assign fifo_intf_1879.wr_en = AESL_inst_myproject.layer3_out_526_U.if_write & AESL_inst_myproject.layer3_out_526_U.if_full_n;
    assign fifo_intf_1879.fifo_rd_block = 0;
    assign fifo_intf_1879.fifo_wr_block = 0;
    assign fifo_intf_1879.finish = finish;
    csv_file_dump fifo_csv_dumper_1879;
    csv_file_dump cstatus_csv_dumper_1879;
    df_fifo_monitor fifo_monitor_1879;
    df_fifo_intf fifo_intf_1880(clock,reset);
    assign fifo_intf_1880.rd_en = AESL_inst_myproject.layer3_out_527_U.if_read & AESL_inst_myproject.layer3_out_527_U.if_empty_n;
    assign fifo_intf_1880.wr_en = AESL_inst_myproject.layer3_out_527_U.if_write & AESL_inst_myproject.layer3_out_527_U.if_full_n;
    assign fifo_intf_1880.fifo_rd_block = 0;
    assign fifo_intf_1880.fifo_wr_block = 0;
    assign fifo_intf_1880.finish = finish;
    csv_file_dump fifo_csv_dumper_1880;
    csv_file_dump cstatus_csv_dumper_1880;
    df_fifo_monitor fifo_monitor_1880;
    df_fifo_intf fifo_intf_1881(clock,reset);
    assign fifo_intf_1881.rd_en = AESL_inst_myproject.layer3_out_528_U.if_read & AESL_inst_myproject.layer3_out_528_U.if_empty_n;
    assign fifo_intf_1881.wr_en = AESL_inst_myproject.layer3_out_528_U.if_write & AESL_inst_myproject.layer3_out_528_U.if_full_n;
    assign fifo_intf_1881.fifo_rd_block = 0;
    assign fifo_intf_1881.fifo_wr_block = 0;
    assign fifo_intf_1881.finish = finish;
    csv_file_dump fifo_csv_dumper_1881;
    csv_file_dump cstatus_csv_dumper_1881;
    df_fifo_monitor fifo_monitor_1881;
    df_fifo_intf fifo_intf_1882(clock,reset);
    assign fifo_intf_1882.rd_en = AESL_inst_myproject.layer3_out_529_U.if_read & AESL_inst_myproject.layer3_out_529_U.if_empty_n;
    assign fifo_intf_1882.wr_en = AESL_inst_myproject.layer3_out_529_U.if_write & AESL_inst_myproject.layer3_out_529_U.if_full_n;
    assign fifo_intf_1882.fifo_rd_block = 0;
    assign fifo_intf_1882.fifo_wr_block = 0;
    assign fifo_intf_1882.finish = finish;
    csv_file_dump fifo_csv_dumper_1882;
    csv_file_dump cstatus_csv_dumper_1882;
    df_fifo_monitor fifo_monitor_1882;
    df_fifo_intf fifo_intf_1883(clock,reset);
    assign fifo_intf_1883.rd_en = AESL_inst_myproject.layer3_out_530_U.if_read & AESL_inst_myproject.layer3_out_530_U.if_empty_n;
    assign fifo_intf_1883.wr_en = AESL_inst_myproject.layer3_out_530_U.if_write & AESL_inst_myproject.layer3_out_530_U.if_full_n;
    assign fifo_intf_1883.fifo_rd_block = 0;
    assign fifo_intf_1883.fifo_wr_block = 0;
    assign fifo_intf_1883.finish = finish;
    csv_file_dump fifo_csv_dumper_1883;
    csv_file_dump cstatus_csv_dumper_1883;
    df_fifo_monitor fifo_monitor_1883;
    df_fifo_intf fifo_intf_1884(clock,reset);
    assign fifo_intf_1884.rd_en = AESL_inst_myproject.layer3_out_531_U.if_read & AESL_inst_myproject.layer3_out_531_U.if_empty_n;
    assign fifo_intf_1884.wr_en = AESL_inst_myproject.layer3_out_531_U.if_write & AESL_inst_myproject.layer3_out_531_U.if_full_n;
    assign fifo_intf_1884.fifo_rd_block = 0;
    assign fifo_intf_1884.fifo_wr_block = 0;
    assign fifo_intf_1884.finish = finish;
    csv_file_dump fifo_csv_dumper_1884;
    csv_file_dump cstatus_csv_dumper_1884;
    df_fifo_monitor fifo_monitor_1884;
    df_fifo_intf fifo_intf_1885(clock,reset);
    assign fifo_intf_1885.rd_en = AESL_inst_myproject.layer3_out_532_U.if_read & AESL_inst_myproject.layer3_out_532_U.if_empty_n;
    assign fifo_intf_1885.wr_en = AESL_inst_myproject.layer3_out_532_U.if_write & AESL_inst_myproject.layer3_out_532_U.if_full_n;
    assign fifo_intf_1885.fifo_rd_block = 0;
    assign fifo_intf_1885.fifo_wr_block = 0;
    assign fifo_intf_1885.finish = finish;
    csv_file_dump fifo_csv_dumper_1885;
    csv_file_dump cstatus_csv_dumper_1885;
    df_fifo_monitor fifo_monitor_1885;
    df_fifo_intf fifo_intf_1886(clock,reset);
    assign fifo_intf_1886.rd_en = AESL_inst_myproject.layer3_out_533_U.if_read & AESL_inst_myproject.layer3_out_533_U.if_empty_n;
    assign fifo_intf_1886.wr_en = AESL_inst_myproject.layer3_out_533_U.if_write & AESL_inst_myproject.layer3_out_533_U.if_full_n;
    assign fifo_intf_1886.fifo_rd_block = 0;
    assign fifo_intf_1886.fifo_wr_block = 0;
    assign fifo_intf_1886.finish = finish;
    csv_file_dump fifo_csv_dumper_1886;
    csv_file_dump cstatus_csv_dumper_1886;
    df_fifo_monitor fifo_monitor_1886;
    df_fifo_intf fifo_intf_1887(clock,reset);
    assign fifo_intf_1887.rd_en = AESL_inst_myproject.layer3_out_534_U.if_read & AESL_inst_myproject.layer3_out_534_U.if_empty_n;
    assign fifo_intf_1887.wr_en = AESL_inst_myproject.layer3_out_534_U.if_write & AESL_inst_myproject.layer3_out_534_U.if_full_n;
    assign fifo_intf_1887.fifo_rd_block = 0;
    assign fifo_intf_1887.fifo_wr_block = 0;
    assign fifo_intf_1887.finish = finish;
    csv_file_dump fifo_csv_dumper_1887;
    csv_file_dump cstatus_csv_dumper_1887;
    df_fifo_monitor fifo_monitor_1887;
    df_fifo_intf fifo_intf_1888(clock,reset);
    assign fifo_intf_1888.rd_en = AESL_inst_myproject.layer3_out_535_U.if_read & AESL_inst_myproject.layer3_out_535_U.if_empty_n;
    assign fifo_intf_1888.wr_en = AESL_inst_myproject.layer3_out_535_U.if_write & AESL_inst_myproject.layer3_out_535_U.if_full_n;
    assign fifo_intf_1888.fifo_rd_block = 0;
    assign fifo_intf_1888.fifo_wr_block = 0;
    assign fifo_intf_1888.finish = finish;
    csv_file_dump fifo_csv_dumper_1888;
    csv_file_dump cstatus_csv_dumper_1888;
    df_fifo_monitor fifo_monitor_1888;
    df_fifo_intf fifo_intf_1889(clock,reset);
    assign fifo_intf_1889.rd_en = AESL_inst_myproject.layer3_out_536_U.if_read & AESL_inst_myproject.layer3_out_536_U.if_empty_n;
    assign fifo_intf_1889.wr_en = AESL_inst_myproject.layer3_out_536_U.if_write & AESL_inst_myproject.layer3_out_536_U.if_full_n;
    assign fifo_intf_1889.fifo_rd_block = 0;
    assign fifo_intf_1889.fifo_wr_block = 0;
    assign fifo_intf_1889.finish = finish;
    csv_file_dump fifo_csv_dumper_1889;
    csv_file_dump cstatus_csv_dumper_1889;
    df_fifo_monitor fifo_monitor_1889;
    df_fifo_intf fifo_intf_1890(clock,reset);
    assign fifo_intf_1890.rd_en = AESL_inst_myproject.layer3_out_537_U.if_read & AESL_inst_myproject.layer3_out_537_U.if_empty_n;
    assign fifo_intf_1890.wr_en = AESL_inst_myproject.layer3_out_537_U.if_write & AESL_inst_myproject.layer3_out_537_U.if_full_n;
    assign fifo_intf_1890.fifo_rd_block = 0;
    assign fifo_intf_1890.fifo_wr_block = 0;
    assign fifo_intf_1890.finish = finish;
    csv_file_dump fifo_csv_dumper_1890;
    csv_file_dump cstatus_csv_dumper_1890;
    df_fifo_monitor fifo_monitor_1890;
    df_fifo_intf fifo_intf_1891(clock,reset);
    assign fifo_intf_1891.rd_en = AESL_inst_myproject.layer3_out_538_U.if_read & AESL_inst_myproject.layer3_out_538_U.if_empty_n;
    assign fifo_intf_1891.wr_en = AESL_inst_myproject.layer3_out_538_U.if_write & AESL_inst_myproject.layer3_out_538_U.if_full_n;
    assign fifo_intf_1891.fifo_rd_block = 0;
    assign fifo_intf_1891.fifo_wr_block = 0;
    assign fifo_intf_1891.finish = finish;
    csv_file_dump fifo_csv_dumper_1891;
    csv_file_dump cstatus_csv_dumper_1891;
    df_fifo_monitor fifo_monitor_1891;
    df_fifo_intf fifo_intf_1892(clock,reset);
    assign fifo_intf_1892.rd_en = AESL_inst_myproject.layer3_out_539_U.if_read & AESL_inst_myproject.layer3_out_539_U.if_empty_n;
    assign fifo_intf_1892.wr_en = AESL_inst_myproject.layer3_out_539_U.if_write & AESL_inst_myproject.layer3_out_539_U.if_full_n;
    assign fifo_intf_1892.fifo_rd_block = 0;
    assign fifo_intf_1892.fifo_wr_block = 0;
    assign fifo_intf_1892.finish = finish;
    csv_file_dump fifo_csv_dumper_1892;
    csv_file_dump cstatus_csv_dumper_1892;
    df_fifo_monitor fifo_monitor_1892;
    df_fifo_intf fifo_intf_1893(clock,reset);
    assign fifo_intf_1893.rd_en = AESL_inst_myproject.layer3_out_540_U.if_read & AESL_inst_myproject.layer3_out_540_U.if_empty_n;
    assign fifo_intf_1893.wr_en = AESL_inst_myproject.layer3_out_540_U.if_write & AESL_inst_myproject.layer3_out_540_U.if_full_n;
    assign fifo_intf_1893.fifo_rd_block = 0;
    assign fifo_intf_1893.fifo_wr_block = 0;
    assign fifo_intf_1893.finish = finish;
    csv_file_dump fifo_csv_dumper_1893;
    csv_file_dump cstatus_csv_dumper_1893;
    df_fifo_monitor fifo_monitor_1893;
    df_fifo_intf fifo_intf_1894(clock,reset);
    assign fifo_intf_1894.rd_en = AESL_inst_myproject.layer3_out_541_U.if_read & AESL_inst_myproject.layer3_out_541_U.if_empty_n;
    assign fifo_intf_1894.wr_en = AESL_inst_myproject.layer3_out_541_U.if_write & AESL_inst_myproject.layer3_out_541_U.if_full_n;
    assign fifo_intf_1894.fifo_rd_block = 0;
    assign fifo_intf_1894.fifo_wr_block = 0;
    assign fifo_intf_1894.finish = finish;
    csv_file_dump fifo_csv_dumper_1894;
    csv_file_dump cstatus_csv_dumper_1894;
    df_fifo_monitor fifo_monitor_1894;
    df_fifo_intf fifo_intf_1895(clock,reset);
    assign fifo_intf_1895.rd_en = AESL_inst_myproject.layer3_out_542_U.if_read & AESL_inst_myproject.layer3_out_542_U.if_empty_n;
    assign fifo_intf_1895.wr_en = AESL_inst_myproject.layer3_out_542_U.if_write & AESL_inst_myproject.layer3_out_542_U.if_full_n;
    assign fifo_intf_1895.fifo_rd_block = 0;
    assign fifo_intf_1895.fifo_wr_block = 0;
    assign fifo_intf_1895.finish = finish;
    csv_file_dump fifo_csv_dumper_1895;
    csv_file_dump cstatus_csv_dumper_1895;
    df_fifo_monitor fifo_monitor_1895;
    df_fifo_intf fifo_intf_1896(clock,reset);
    assign fifo_intf_1896.rd_en = AESL_inst_myproject.layer3_out_543_U.if_read & AESL_inst_myproject.layer3_out_543_U.if_empty_n;
    assign fifo_intf_1896.wr_en = AESL_inst_myproject.layer3_out_543_U.if_write & AESL_inst_myproject.layer3_out_543_U.if_full_n;
    assign fifo_intf_1896.fifo_rd_block = 0;
    assign fifo_intf_1896.fifo_wr_block = 0;
    assign fifo_intf_1896.finish = finish;
    csv_file_dump fifo_csv_dumper_1896;
    csv_file_dump cstatus_csv_dumper_1896;
    df_fifo_monitor fifo_monitor_1896;
    df_fifo_intf fifo_intf_1897(clock,reset);
    assign fifo_intf_1897.rd_en = AESL_inst_myproject.layer3_out_544_U.if_read & AESL_inst_myproject.layer3_out_544_U.if_empty_n;
    assign fifo_intf_1897.wr_en = AESL_inst_myproject.layer3_out_544_U.if_write & AESL_inst_myproject.layer3_out_544_U.if_full_n;
    assign fifo_intf_1897.fifo_rd_block = 0;
    assign fifo_intf_1897.fifo_wr_block = 0;
    assign fifo_intf_1897.finish = finish;
    csv_file_dump fifo_csv_dumper_1897;
    csv_file_dump cstatus_csv_dumper_1897;
    df_fifo_monitor fifo_monitor_1897;
    df_fifo_intf fifo_intf_1898(clock,reset);
    assign fifo_intf_1898.rd_en = AESL_inst_myproject.layer3_out_545_U.if_read & AESL_inst_myproject.layer3_out_545_U.if_empty_n;
    assign fifo_intf_1898.wr_en = AESL_inst_myproject.layer3_out_545_U.if_write & AESL_inst_myproject.layer3_out_545_U.if_full_n;
    assign fifo_intf_1898.fifo_rd_block = 0;
    assign fifo_intf_1898.fifo_wr_block = 0;
    assign fifo_intf_1898.finish = finish;
    csv_file_dump fifo_csv_dumper_1898;
    csv_file_dump cstatus_csv_dumper_1898;
    df_fifo_monitor fifo_monitor_1898;
    df_fifo_intf fifo_intf_1899(clock,reset);
    assign fifo_intf_1899.rd_en = AESL_inst_myproject.layer3_out_546_U.if_read & AESL_inst_myproject.layer3_out_546_U.if_empty_n;
    assign fifo_intf_1899.wr_en = AESL_inst_myproject.layer3_out_546_U.if_write & AESL_inst_myproject.layer3_out_546_U.if_full_n;
    assign fifo_intf_1899.fifo_rd_block = 0;
    assign fifo_intf_1899.fifo_wr_block = 0;
    assign fifo_intf_1899.finish = finish;
    csv_file_dump fifo_csv_dumper_1899;
    csv_file_dump cstatus_csv_dumper_1899;
    df_fifo_monitor fifo_monitor_1899;
    df_fifo_intf fifo_intf_1900(clock,reset);
    assign fifo_intf_1900.rd_en = AESL_inst_myproject.layer3_out_547_U.if_read & AESL_inst_myproject.layer3_out_547_U.if_empty_n;
    assign fifo_intf_1900.wr_en = AESL_inst_myproject.layer3_out_547_U.if_write & AESL_inst_myproject.layer3_out_547_U.if_full_n;
    assign fifo_intf_1900.fifo_rd_block = 0;
    assign fifo_intf_1900.fifo_wr_block = 0;
    assign fifo_intf_1900.finish = finish;
    csv_file_dump fifo_csv_dumper_1900;
    csv_file_dump cstatus_csv_dumper_1900;
    df_fifo_monitor fifo_monitor_1900;
    df_fifo_intf fifo_intf_1901(clock,reset);
    assign fifo_intf_1901.rd_en = AESL_inst_myproject.layer3_out_548_U.if_read & AESL_inst_myproject.layer3_out_548_U.if_empty_n;
    assign fifo_intf_1901.wr_en = AESL_inst_myproject.layer3_out_548_U.if_write & AESL_inst_myproject.layer3_out_548_U.if_full_n;
    assign fifo_intf_1901.fifo_rd_block = 0;
    assign fifo_intf_1901.fifo_wr_block = 0;
    assign fifo_intf_1901.finish = finish;
    csv_file_dump fifo_csv_dumper_1901;
    csv_file_dump cstatus_csv_dumper_1901;
    df_fifo_monitor fifo_monitor_1901;
    df_fifo_intf fifo_intf_1902(clock,reset);
    assign fifo_intf_1902.rd_en = AESL_inst_myproject.layer3_out_549_U.if_read & AESL_inst_myproject.layer3_out_549_U.if_empty_n;
    assign fifo_intf_1902.wr_en = AESL_inst_myproject.layer3_out_549_U.if_write & AESL_inst_myproject.layer3_out_549_U.if_full_n;
    assign fifo_intf_1902.fifo_rd_block = 0;
    assign fifo_intf_1902.fifo_wr_block = 0;
    assign fifo_intf_1902.finish = finish;
    csv_file_dump fifo_csv_dumper_1902;
    csv_file_dump cstatus_csv_dumper_1902;
    df_fifo_monitor fifo_monitor_1902;
    df_fifo_intf fifo_intf_1903(clock,reset);
    assign fifo_intf_1903.rd_en = AESL_inst_myproject.layer3_out_550_U.if_read & AESL_inst_myproject.layer3_out_550_U.if_empty_n;
    assign fifo_intf_1903.wr_en = AESL_inst_myproject.layer3_out_550_U.if_write & AESL_inst_myproject.layer3_out_550_U.if_full_n;
    assign fifo_intf_1903.fifo_rd_block = 0;
    assign fifo_intf_1903.fifo_wr_block = 0;
    assign fifo_intf_1903.finish = finish;
    csv_file_dump fifo_csv_dumper_1903;
    csv_file_dump cstatus_csv_dumper_1903;
    df_fifo_monitor fifo_monitor_1903;
    df_fifo_intf fifo_intf_1904(clock,reset);
    assign fifo_intf_1904.rd_en = AESL_inst_myproject.layer3_out_551_U.if_read & AESL_inst_myproject.layer3_out_551_U.if_empty_n;
    assign fifo_intf_1904.wr_en = AESL_inst_myproject.layer3_out_551_U.if_write & AESL_inst_myproject.layer3_out_551_U.if_full_n;
    assign fifo_intf_1904.fifo_rd_block = 0;
    assign fifo_intf_1904.fifo_wr_block = 0;
    assign fifo_intf_1904.finish = finish;
    csv_file_dump fifo_csv_dumper_1904;
    csv_file_dump cstatus_csv_dumper_1904;
    df_fifo_monitor fifo_monitor_1904;
    df_fifo_intf fifo_intf_1905(clock,reset);
    assign fifo_intf_1905.rd_en = AESL_inst_myproject.layer3_out_552_U.if_read & AESL_inst_myproject.layer3_out_552_U.if_empty_n;
    assign fifo_intf_1905.wr_en = AESL_inst_myproject.layer3_out_552_U.if_write & AESL_inst_myproject.layer3_out_552_U.if_full_n;
    assign fifo_intf_1905.fifo_rd_block = 0;
    assign fifo_intf_1905.fifo_wr_block = 0;
    assign fifo_intf_1905.finish = finish;
    csv_file_dump fifo_csv_dumper_1905;
    csv_file_dump cstatus_csv_dumper_1905;
    df_fifo_monitor fifo_monitor_1905;
    df_fifo_intf fifo_intf_1906(clock,reset);
    assign fifo_intf_1906.rd_en = AESL_inst_myproject.layer3_out_553_U.if_read & AESL_inst_myproject.layer3_out_553_U.if_empty_n;
    assign fifo_intf_1906.wr_en = AESL_inst_myproject.layer3_out_553_U.if_write & AESL_inst_myproject.layer3_out_553_U.if_full_n;
    assign fifo_intf_1906.fifo_rd_block = 0;
    assign fifo_intf_1906.fifo_wr_block = 0;
    assign fifo_intf_1906.finish = finish;
    csv_file_dump fifo_csv_dumper_1906;
    csv_file_dump cstatus_csv_dumper_1906;
    df_fifo_monitor fifo_monitor_1906;
    df_fifo_intf fifo_intf_1907(clock,reset);
    assign fifo_intf_1907.rd_en = AESL_inst_myproject.layer3_out_554_U.if_read & AESL_inst_myproject.layer3_out_554_U.if_empty_n;
    assign fifo_intf_1907.wr_en = AESL_inst_myproject.layer3_out_554_U.if_write & AESL_inst_myproject.layer3_out_554_U.if_full_n;
    assign fifo_intf_1907.fifo_rd_block = 0;
    assign fifo_intf_1907.fifo_wr_block = 0;
    assign fifo_intf_1907.finish = finish;
    csv_file_dump fifo_csv_dumper_1907;
    csv_file_dump cstatus_csv_dumper_1907;
    df_fifo_monitor fifo_monitor_1907;
    df_fifo_intf fifo_intf_1908(clock,reset);
    assign fifo_intf_1908.rd_en = AESL_inst_myproject.layer3_out_555_U.if_read & AESL_inst_myproject.layer3_out_555_U.if_empty_n;
    assign fifo_intf_1908.wr_en = AESL_inst_myproject.layer3_out_555_U.if_write & AESL_inst_myproject.layer3_out_555_U.if_full_n;
    assign fifo_intf_1908.fifo_rd_block = 0;
    assign fifo_intf_1908.fifo_wr_block = 0;
    assign fifo_intf_1908.finish = finish;
    csv_file_dump fifo_csv_dumper_1908;
    csv_file_dump cstatus_csv_dumper_1908;
    df_fifo_monitor fifo_monitor_1908;
    df_fifo_intf fifo_intf_1909(clock,reset);
    assign fifo_intf_1909.rd_en = AESL_inst_myproject.layer3_out_556_U.if_read & AESL_inst_myproject.layer3_out_556_U.if_empty_n;
    assign fifo_intf_1909.wr_en = AESL_inst_myproject.layer3_out_556_U.if_write & AESL_inst_myproject.layer3_out_556_U.if_full_n;
    assign fifo_intf_1909.fifo_rd_block = 0;
    assign fifo_intf_1909.fifo_wr_block = 0;
    assign fifo_intf_1909.finish = finish;
    csv_file_dump fifo_csv_dumper_1909;
    csv_file_dump cstatus_csv_dumper_1909;
    df_fifo_monitor fifo_monitor_1909;
    df_fifo_intf fifo_intf_1910(clock,reset);
    assign fifo_intf_1910.rd_en = AESL_inst_myproject.layer3_out_557_U.if_read & AESL_inst_myproject.layer3_out_557_U.if_empty_n;
    assign fifo_intf_1910.wr_en = AESL_inst_myproject.layer3_out_557_U.if_write & AESL_inst_myproject.layer3_out_557_U.if_full_n;
    assign fifo_intf_1910.fifo_rd_block = 0;
    assign fifo_intf_1910.fifo_wr_block = 0;
    assign fifo_intf_1910.finish = finish;
    csv_file_dump fifo_csv_dumper_1910;
    csv_file_dump cstatus_csv_dumper_1910;
    df_fifo_monitor fifo_monitor_1910;
    df_fifo_intf fifo_intf_1911(clock,reset);
    assign fifo_intf_1911.rd_en = AESL_inst_myproject.layer3_out_558_U.if_read & AESL_inst_myproject.layer3_out_558_U.if_empty_n;
    assign fifo_intf_1911.wr_en = AESL_inst_myproject.layer3_out_558_U.if_write & AESL_inst_myproject.layer3_out_558_U.if_full_n;
    assign fifo_intf_1911.fifo_rd_block = 0;
    assign fifo_intf_1911.fifo_wr_block = 0;
    assign fifo_intf_1911.finish = finish;
    csv_file_dump fifo_csv_dumper_1911;
    csv_file_dump cstatus_csv_dumper_1911;
    df_fifo_monitor fifo_monitor_1911;
    df_fifo_intf fifo_intf_1912(clock,reset);
    assign fifo_intf_1912.rd_en = AESL_inst_myproject.layer3_out_559_U.if_read & AESL_inst_myproject.layer3_out_559_U.if_empty_n;
    assign fifo_intf_1912.wr_en = AESL_inst_myproject.layer3_out_559_U.if_write & AESL_inst_myproject.layer3_out_559_U.if_full_n;
    assign fifo_intf_1912.fifo_rd_block = 0;
    assign fifo_intf_1912.fifo_wr_block = 0;
    assign fifo_intf_1912.finish = finish;
    csv_file_dump fifo_csv_dumper_1912;
    csv_file_dump cstatus_csv_dumper_1912;
    df_fifo_monitor fifo_monitor_1912;
    df_fifo_intf fifo_intf_1913(clock,reset);
    assign fifo_intf_1913.rd_en = AESL_inst_myproject.layer3_out_560_U.if_read & AESL_inst_myproject.layer3_out_560_U.if_empty_n;
    assign fifo_intf_1913.wr_en = AESL_inst_myproject.layer3_out_560_U.if_write & AESL_inst_myproject.layer3_out_560_U.if_full_n;
    assign fifo_intf_1913.fifo_rd_block = 0;
    assign fifo_intf_1913.fifo_wr_block = 0;
    assign fifo_intf_1913.finish = finish;
    csv_file_dump fifo_csv_dumper_1913;
    csv_file_dump cstatus_csv_dumper_1913;
    df_fifo_monitor fifo_monitor_1913;
    df_fifo_intf fifo_intf_1914(clock,reset);
    assign fifo_intf_1914.rd_en = AESL_inst_myproject.layer3_out_561_U.if_read & AESL_inst_myproject.layer3_out_561_U.if_empty_n;
    assign fifo_intf_1914.wr_en = AESL_inst_myproject.layer3_out_561_U.if_write & AESL_inst_myproject.layer3_out_561_U.if_full_n;
    assign fifo_intf_1914.fifo_rd_block = 0;
    assign fifo_intf_1914.fifo_wr_block = 0;
    assign fifo_intf_1914.finish = finish;
    csv_file_dump fifo_csv_dumper_1914;
    csv_file_dump cstatus_csv_dumper_1914;
    df_fifo_monitor fifo_monitor_1914;
    df_fifo_intf fifo_intf_1915(clock,reset);
    assign fifo_intf_1915.rd_en = AESL_inst_myproject.layer3_out_562_U.if_read & AESL_inst_myproject.layer3_out_562_U.if_empty_n;
    assign fifo_intf_1915.wr_en = AESL_inst_myproject.layer3_out_562_U.if_write & AESL_inst_myproject.layer3_out_562_U.if_full_n;
    assign fifo_intf_1915.fifo_rd_block = 0;
    assign fifo_intf_1915.fifo_wr_block = 0;
    assign fifo_intf_1915.finish = finish;
    csv_file_dump fifo_csv_dumper_1915;
    csv_file_dump cstatus_csv_dumper_1915;
    df_fifo_monitor fifo_monitor_1915;
    df_fifo_intf fifo_intf_1916(clock,reset);
    assign fifo_intf_1916.rd_en = AESL_inst_myproject.layer3_out_563_U.if_read & AESL_inst_myproject.layer3_out_563_U.if_empty_n;
    assign fifo_intf_1916.wr_en = AESL_inst_myproject.layer3_out_563_U.if_write & AESL_inst_myproject.layer3_out_563_U.if_full_n;
    assign fifo_intf_1916.fifo_rd_block = 0;
    assign fifo_intf_1916.fifo_wr_block = 0;
    assign fifo_intf_1916.finish = finish;
    csv_file_dump fifo_csv_dumper_1916;
    csv_file_dump cstatus_csv_dumper_1916;
    df_fifo_monitor fifo_monitor_1916;
    df_fifo_intf fifo_intf_1917(clock,reset);
    assign fifo_intf_1917.rd_en = AESL_inst_myproject.layer3_out_564_U.if_read & AESL_inst_myproject.layer3_out_564_U.if_empty_n;
    assign fifo_intf_1917.wr_en = AESL_inst_myproject.layer3_out_564_U.if_write & AESL_inst_myproject.layer3_out_564_U.if_full_n;
    assign fifo_intf_1917.fifo_rd_block = 0;
    assign fifo_intf_1917.fifo_wr_block = 0;
    assign fifo_intf_1917.finish = finish;
    csv_file_dump fifo_csv_dumper_1917;
    csv_file_dump cstatus_csv_dumper_1917;
    df_fifo_monitor fifo_monitor_1917;
    df_fifo_intf fifo_intf_1918(clock,reset);
    assign fifo_intf_1918.rd_en = AESL_inst_myproject.layer3_out_565_U.if_read & AESL_inst_myproject.layer3_out_565_U.if_empty_n;
    assign fifo_intf_1918.wr_en = AESL_inst_myproject.layer3_out_565_U.if_write & AESL_inst_myproject.layer3_out_565_U.if_full_n;
    assign fifo_intf_1918.fifo_rd_block = 0;
    assign fifo_intf_1918.fifo_wr_block = 0;
    assign fifo_intf_1918.finish = finish;
    csv_file_dump fifo_csv_dumper_1918;
    csv_file_dump cstatus_csv_dumper_1918;
    df_fifo_monitor fifo_monitor_1918;
    df_fifo_intf fifo_intf_1919(clock,reset);
    assign fifo_intf_1919.rd_en = AESL_inst_myproject.layer3_out_566_U.if_read & AESL_inst_myproject.layer3_out_566_U.if_empty_n;
    assign fifo_intf_1919.wr_en = AESL_inst_myproject.layer3_out_566_U.if_write & AESL_inst_myproject.layer3_out_566_U.if_full_n;
    assign fifo_intf_1919.fifo_rd_block = 0;
    assign fifo_intf_1919.fifo_wr_block = 0;
    assign fifo_intf_1919.finish = finish;
    csv_file_dump fifo_csv_dumper_1919;
    csv_file_dump cstatus_csv_dumper_1919;
    df_fifo_monitor fifo_monitor_1919;
    df_fifo_intf fifo_intf_1920(clock,reset);
    assign fifo_intf_1920.rd_en = AESL_inst_myproject.layer3_out_567_U.if_read & AESL_inst_myproject.layer3_out_567_U.if_empty_n;
    assign fifo_intf_1920.wr_en = AESL_inst_myproject.layer3_out_567_U.if_write & AESL_inst_myproject.layer3_out_567_U.if_full_n;
    assign fifo_intf_1920.fifo_rd_block = 0;
    assign fifo_intf_1920.fifo_wr_block = 0;
    assign fifo_intf_1920.finish = finish;
    csv_file_dump fifo_csv_dumper_1920;
    csv_file_dump cstatus_csv_dumper_1920;
    df_fifo_monitor fifo_monitor_1920;
    df_fifo_intf fifo_intf_1921(clock,reset);
    assign fifo_intf_1921.rd_en = AESL_inst_myproject.layer3_out_568_U.if_read & AESL_inst_myproject.layer3_out_568_U.if_empty_n;
    assign fifo_intf_1921.wr_en = AESL_inst_myproject.layer3_out_568_U.if_write & AESL_inst_myproject.layer3_out_568_U.if_full_n;
    assign fifo_intf_1921.fifo_rd_block = 0;
    assign fifo_intf_1921.fifo_wr_block = 0;
    assign fifo_intf_1921.finish = finish;
    csv_file_dump fifo_csv_dumper_1921;
    csv_file_dump cstatus_csv_dumper_1921;
    df_fifo_monitor fifo_monitor_1921;
    df_fifo_intf fifo_intf_1922(clock,reset);
    assign fifo_intf_1922.rd_en = AESL_inst_myproject.layer3_out_569_U.if_read & AESL_inst_myproject.layer3_out_569_U.if_empty_n;
    assign fifo_intf_1922.wr_en = AESL_inst_myproject.layer3_out_569_U.if_write & AESL_inst_myproject.layer3_out_569_U.if_full_n;
    assign fifo_intf_1922.fifo_rd_block = 0;
    assign fifo_intf_1922.fifo_wr_block = 0;
    assign fifo_intf_1922.finish = finish;
    csv_file_dump fifo_csv_dumper_1922;
    csv_file_dump cstatus_csv_dumper_1922;
    df_fifo_monitor fifo_monitor_1922;
    df_fifo_intf fifo_intf_1923(clock,reset);
    assign fifo_intf_1923.rd_en = AESL_inst_myproject.layer3_out_570_U.if_read & AESL_inst_myproject.layer3_out_570_U.if_empty_n;
    assign fifo_intf_1923.wr_en = AESL_inst_myproject.layer3_out_570_U.if_write & AESL_inst_myproject.layer3_out_570_U.if_full_n;
    assign fifo_intf_1923.fifo_rd_block = 0;
    assign fifo_intf_1923.fifo_wr_block = 0;
    assign fifo_intf_1923.finish = finish;
    csv_file_dump fifo_csv_dumper_1923;
    csv_file_dump cstatus_csv_dumper_1923;
    df_fifo_monitor fifo_monitor_1923;
    df_fifo_intf fifo_intf_1924(clock,reset);
    assign fifo_intf_1924.rd_en = AESL_inst_myproject.layer3_out_571_U.if_read & AESL_inst_myproject.layer3_out_571_U.if_empty_n;
    assign fifo_intf_1924.wr_en = AESL_inst_myproject.layer3_out_571_U.if_write & AESL_inst_myproject.layer3_out_571_U.if_full_n;
    assign fifo_intf_1924.fifo_rd_block = 0;
    assign fifo_intf_1924.fifo_wr_block = 0;
    assign fifo_intf_1924.finish = finish;
    csv_file_dump fifo_csv_dumper_1924;
    csv_file_dump cstatus_csv_dumper_1924;
    df_fifo_monitor fifo_monitor_1924;
    df_fifo_intf fifo_intf_1925(clock,reset);
    assign fifo_intf_1925.rd_en = AESL_inst_myproject.layer3_out_572_U.if_read & AESL_inst_myproject.layer3_out_572_U.if_empty_n;
    assign fifo_intf_1925.wr_en = AESL_inst_myproject.layer3_out_572_U.if_write & AESL_inst_myproject.layer3_out_572_U.if_full_n;
    assign fifo_intf_1925.fifo_rd_block = 0;
    assign fifo_intf_1925.fifo_wr_block = 0;
    assign fifo_intf_1925.finish = finish;
    csv_file_dump fifo_csv_dumper_1925;
    csv_file_dump cstatus_csv_dumper_1925;
    df_fifo_monitor fifo_monitor_1925;
    df_fifo_intf fifo_intf_1926(clock,reset);
    assign fifo_intf_1926.rd_en = AESL_inst_myproject.layer3_out_573_U.if_read & AESL_inst_myproject.layer3_out_573_U.if_empty_n;
    assign fifo_intf_1926.wr_en = AESL_inst_myproject.layer3_out_573_U.if_write & AESL_inst_myproject.layer3_out_573_U.if_full_n;
    assign fifo_intf_1926.fifo_rd_block = 0;
    assign fifo_intf_1926.fifo_wr_block = 0;
    assign fifo_intf_1926.finish = finish;
    csv_file_dump fifo_csv_dumper_1926;
    csv_file_dump cstatus_csv_dumper_1926;
    df_fifo_monitor fifo_monitor_1926;
    df_fifo_intf fifo_intf_1927(clock,reset);
    assign fifo_intf_1927.rd_en = AESL_inst_myproject.layer3_out_574_U.if_read & AESL_inst_myproject.layer3_out_574_U.if_empty_n;
    assign fifo_intf_1927.wr_en = AESL_inst_myproject.layer3_out_574_U.if_write & AESL_inst_myproject.layer3_out_574_U.if_full_n;
    assign fifo_intf_1927.fifo_rd_block = 0;
    assign fifo_intf_1927.fifo_wr_block = 0;
    assign fifo_intf_1927.finish = finish;
    csv_file_dump fifo_csv_dumper_1927;
    csv_file_dump cstatus_csv_dumper_1927;
    df_fifo_monitor fifo_monitor_1927;
    df_fifo_intf fifo_intf_1928(clock,reset);
    assign fifo_intf_1928.rd_en = AESL_inst_myproject.layer3_out_575_U.if_read & AESL_inst_myproject.layer3_out_575_U.if_empty_n;
    assign fifo_intf_1928.wr_en = AESL_inst_myproject.layer3_out_575_U.if_write & AESL_inst_myproject.layer3_out_575_U.if_full_n;
    assign fifo_intf_1928.fifo_rd_block = 0;
    assign fifo_intf_1928.fifo_wr_block = 0;
    assign fifo_intf_1928.finish = finish;
    csv_file_dump fifo_csv_dumper_1928;
    csv_file_dump cstatus_csv_dumper_1928;
    df_fifo_monitor fifo_monitor_1928;
    df_fifo_intf fifo_intf_1929(clock,reset);
    assign fifo_intf_1929.rd_en = AESL_inst_myproject.layer3_out_576_U.if_read & AESL_inst_myproject.layer3_out_576_U.if_empty_n;
    assign fifo_intf_1929.wr_en = AESL_inst_myproject.layer3_out_576_U.if_write & AESL_inst_myproject.layer3_out_576_U.if_full_n;
    assign fifo_intf_1929.fifo_rd_block = 0;
    assign fifo_intf_1929.fifo_wr_block = 0;
    assign fifo_intf_1929.finish = finish;
    csv_file_dump fifo_csv_dumper_1929;
    csv_file_dump cstatus_csv_dumper_1929;
    df_fifo_monitor fifo_monitor_1929;
    df_fifo_intf fifo_intf_1930(clock,reset);
    assign fifo_intf_1930.rd_en = AESL_inst_myproject.layer3_out_577_U.if_read & AESL_inst_myproject.layer3_out_577_U.if_empty_n;
    assign fifo_intf_1930.wr_en = AESL_inst_myproject.layer3_out_577_U.if_write & AESL_inst_myproject.layer3_out_577_U.if_full_n;
    assign fifo_intf_1930.fifo_rd_block = 0;
    assign fifo_intf_1930.fifo_wr_block = 0;
    assign fifo_intf_1930.finish = finish;
    csv_file_dump fifo_csv_dumper_1930;
    csv_file_dump cstatus_csv_dumper_1930;
    df_fifo_monitor fifo_monitor_1930;
    df_fifo_intf fifo_intf_1931(clock,reset);
    assign fifo_intf_1931.rd_en = AESL_inst_myproject.layer3_out_578_U.if_read & AESL_inst_myproject.layer3_out_578_U.if_empty_n;
    assign fifo_intf_1931.wr_en = AESL_inst_myproject.layer3_out_578_U.if_write & AESL_inst_myproject.layer3_out_578_U.if_full_n;
    assign fifo_intf_1931.fifo_rd_block = 0;
    assign fifo_intf_1931.fifo_wr_block = 0;
    assign fifo_intf_1931.finish = finish;
    csv_file_dump fifo_csv_dumper_1931;
    csv_file_dump cstatus_csv_dumper_1931;
    df_fifo_monitor fifo_monitor_1931;
    df_fifo_intf fifo_intf_1932(clock,reset);
    assign fifo_intf_1932.rd_en = AESL_inst_myproject.layer3_out_579_U.if_read & AESL_inst_myproject.layer3_out_579_U.if_empty_n;
    assign fifo_intf_1932.wr_en = AESL_inst_myproject.layer3_out_579_U.if_write & AESL_inst_myproject.layer3_out_579_U.if_full_n;
    assign fifo_intf_1932.fifo_rd_block = 0;
    assign fifo_intf_1932.fifo_wr_block = 0;
    assign fifo_intf_1932.finish = finish;
    csv_file_dump fifo_csv_dumper_1932;
    csv_file_dump cstatus_csv_dumper_1932;
    df_fifo_monitor fifo_monitor_1932;
    df_fifo_intf fifo_intf_1933(clock,reset);
    assign fifo_intf_1933.rd_en = AESL_inst_myproject.layer3_out_580_U.if_read & AESL_inst_myproject.layer3_out_580_U.if_empty_n;
    assign fifo_intf_1933.wr_en = AESL_inst_myproject.layer3_out_580_U.if_write & AESL_inst_myproject.layer3_out_580_U.if_full_n;
    assign fifo_intf_1933.fifo_rd_block = 0;
    assign fifo_intf_1933.fifo_wr_block = 0;
    assign fifo_intf_1933.finish = finish;
    csv_file_dump fifo_csv_dumper_1933;
    csv_file_dump cstatus_csv_dumper_1933;
    df_fifo_monitor fifo_monitor_1933;
    df_fifo_intf fifo_intf_1934(clock,reset);
    assign fifo_intf_1934.rd_en = AESL_inst_myproject.layer3_out_581_U.if_read & AESL_inst_myproject.layer3_out_581_U.if_empty_n;
    assign fifo_intf_1934.wr_en = AESL_inst_myproject.layer3_out_581_U.if_write & AESL_inst_myproject.layer3_out_581_U.if_full_n;
    assign fifo_intf_1934.fifo_rd_block = 0;
    assign fifo_intf_1934.fifo_wr_block = 0;
    assign fifo_intf_1934.finish = finish;
    csv_file_dump fifo_csv_dumper_1934;
    csv_file_dump cstatus_csv_dumper_1934;
    df_fifo_monitor fifo_monitor_1934;
    df_fifo_intf fifo_intf_1935(clock,reset);
    assign fifo_intf_1935.rd_en = AESL_inst_myproject.layer3_out_582_U.if_read & AESL_inst_myproject.layer3_out_582_U.if_empty_n;
    assign fifo_intf_1935.wr_en = AESL_inst_myproject.layer3_out_582_U.if_write & AESL_inst_myproject.layer3_out_582_U.if_full_n;
    assign fifo_intf_1935.fifo_rd_block = 0;
    assign fifo_intf_1935.fifo_wr_block = 0;
    assign fifo_intf_1935.finish = finish;
    csv_file_dump fifo_csv_dumper_1935;
    csv_file_dump cstatus_csv_dumper_1935;
    df_fifo_monitor fifo_monitor_1935;
    df_fifo_intf fifo_intf_1936(clock,reset);
    assign fifo_intf_1936.rd_en = AESL_inst_myproject.layer3_out_583_U.if_read & AESL_inst_myproject.layer3_out_583_U.if_empty_n;
    assign fifo_intf_1936.wr_en = AESL_inst_myproject.layer3_out_583_U.if_write & AESL_inst_myproject.layer3_out_583_U.if_full_n;
    assign fifo_intf_1936.fifo_rd_block = 0;
    assign fifo_intf_1936.fifo_wr_block = 0;
    assign fifo_intf_1936.finish = finish;
    csv_file_dump fifo_csv_dumper_1936;
    csv_file_dump cstatus_csv_dumper_1936;
    df_fifo_monitor fifo_monitor_1936;
    df_fifo_intf fifo_intf_1937(clock,reset);
    assign fifo_intf_1937.rd_en = AESL_inst_myproject.layer3_out_584_U.if_read & AESL_inst_myproject.layer3_out_584_U.if_empty_n;
    assign fifo_intf_1937.wr_en = AESL_inst_myproject.layer3_out_584_U.if_write & AESL_inst_myproject.layer3_out_584_U.if_full_n;
    assign fifo_intf_1937.fifo_rd_block = 0;
    assign fifo_intf_1937.fifo_wr_block = 0;
    assign fifo_intf_1937.finish = finish;
    csv_file_dump fifo_csv_dumper_1937;
    csv_file_dump cstatus_csv_dumper_1937;
    df_fifo_monitor fifo_monitor_1937;
    df_fifo_intf fifo_intf_1938(clock,reset);
    assign fifo_intf_1938.rd_en = AESL_inst_myproject.layer3_out_585_U.if_read & AESL_inst_myproject.layer3_out_585_U.if_empty_n;
    assign fifo_intf_1938.wr_en = AESL_inst_myproject.layer3_out_585_U.if_write & AESL_inst_myproject.layer3_out_585_U.if_full_n;
    assign fifo_intf_1938.fifo_rd_block = 0;
    assign fifo_intf_1938.fifo_wr_block = 0;
    assign fifo_intf_1938.finish = finish;
    csv_file_dump fifo_csv_dumper_1938;
    csv_file_dump cstatus_csv_dumper_1938;
    df_fifo_monitor fifo_monitor_1938;
    df_fifo_intf fifo_intf_1939(clock,reset);
    assign fifo_intf_1939.rd_en = AESL_inst_myproject.layer3_out_586_U.if_read & AESL_inst_myproject.layer3_out_586_U.if_empty_n;
    assign fifo_intf_1939.wr_en = AESL_inst_myproject.layer3_out_586_U.if_write & AESL_inst_myproject.layer3_out_586_U.if_full_n;
    assign fifo_intf_1939.fifo_rd_block = 0;
    assign fifo_intf_1939.fifo_wr_block = 0;
    assign fifo_intf_1939.finish = finish;
    csv_file_dump fifo_csv_dumper_1939;
    csv_file_dump cstatus_csv_dumper_1939;
    df_fifo_monitor fifo_monitor_1939;
    df_fifo_intf fifo_intf_1940(clock,reset);
    assign fifo_intf_1940.rd_en = AESL_inst_myproject.layer3_out_587_U.if_read & AESL_inst_myproject.layer3_out_587_U.if_empty_n;
    assign fifo_intf_1940.wr_en = AESL_inst_myproject.layer3_out_587_U.if_write & AESL_inst_myproject.layer3_out_587_U.if_full_n;
    assign fifo_intf_1940.fifo_rd_block = 0;
    assign fifo_intf_1940.fifo_wr_block = 0;
    assign fifo_intf_1940.finish = finish;
    csv_file_dump fifo_csv_dumper_1940;
    csv_file_dump cstatus_csv_dumper_1940;
    df_fifo_monitor fifo_monitor_1940;
    df_fifo_intf fifo_intf_1941(clock,reset);
    assign fifo_intf_1941.rd_en = AESL_inst_myproject.layer3_out_588_U.if_read & AESL_inst_myproject.layer3_out_588_U.if_empty_n;
    assign fifo_intf_1941.wr_en = AESL_inst_myproject.layer3_out_588_U.if_write & AESL_inst_myproject.layer3_out_588_U.if_full_n;
    assign fifo_intf_1941.fifo_rd_block = 0;
    assign fifo_intf_1941.fifo_wr_block = 0;
    assign fifo_intf_1941.finish = finish;
    csv_file_dump fifo_csv_dumper_1941;
    csv_file_dump cstatus_csv_dumper_1941;
    df_fifo_monitor fifo_monitor_1941;
    df_fifo_intf fifo_intf_1942(clock,reset);
    assign fifo_intf_1942.rd_en = AESL_inst_myproject.layer3_out_589_U.if_read & AESL_inst_myproject.layer3_out_589_U.if_empty_n;
    assign fifo_intf_1942.wr_en = AESL_inst_myproject.layer3_out_589_U.if_write & AESL_inst_myproject.layer3_out_589_U.if_full_n;
    assign fifo_intf_1942.fifo_rd_block = 0;
    assign fifo_intf_1942.fifo_wr_block = 0;
    assign fifo_intf_1942.finish = finish;
    csv_file_dump fifo_csv_dumper_1942;
    csv_file_dump cstatus_csv_dumper_1942;
    df_fifo_monitor fifo_monitor_1942;
    df_fifo_intf fifo_intf_1943(clock,reset);
    assign fifo_intf_1943.rd_en = AESL_inst_myproject.layer3_out_590_U.if_read & AESL_inst_myproject.layer3_out_590_U.if_empty_n;
    assign fifo_intf_1943.wr_en = AESL_inst_myproject.layer3_out_590_U.if_write & AESL_inst_myproject.layer3_out_590_U.if_full_n;
    assign fifo_intf_1943.fifo_rd_block = 0;
    assign fifo_intf_1943.fifo_wr_block = 0;
    assign fifo_intf_1943.finish = finish;
    csv_file_dump fifo_csv_dumper_1943;
    csv_file_dump cstatus_csv_dumper_1943;
    df_fifo_monitor fifo_monitor_1943;
    df_fifo_intf fifo_intf_1944(clock,reset);
    assign fifo_intf_1944.rd_en = AESL_inst_myproject.layer3_out_591_U.if_read & AESL_inst_myproject.layer3_out_591_U.if_empty_n;
    assign fifo_intf_1944.wr_en = AESL_inst_myproject.layer3_out_591_U.if_write & AESL_inst_myproject.layer3_out_591_U.if_full_n;
    assign fifo_intf_1944.fifo_rd_block = 0;
    assign fifo_intf_1944.fifo_wr_block = 0;
    assign fifo_intf_1944.finish = finish;
    csv_file_dump fifo_csv_dumper_1944;
    csv_file_dump cstatus_csv_dumper_1944;
    df_fifo_monitor fifo_monitor_1944;
    df_fifo_intf fifo_intf_1945(clock,reset);
    assign fifo_intf_1945.rd_en = AESL_inst_myproject.layer3_out_592_U.if_read & AESL_inst_myproject.layer3_out_592_U.if_empty_n;
    assign fifo_intf_1945.wr_en = AESL_inst_myproject.layer3_out_592_U.if_write & AESL_inst_myproject.layer3_out_592_U.if_full_n;
    assign fifo_intf_1945.fifo_rd_block = 0;
    assign fifo_intf_1945.fifo_wr_block = 0;
    assign fifo_intf_1945.finish = finish;
    csv_file_dump fifo_csv_dumper_1945;
    csv_file_dump cstatus_csv_dumper_1945;
    df_fifo_monitor fifo_monitor_1945;
    df_fifo_intf fifo_intf_1946(clock,reset);
    assign fifo_intf_1946.rd_en = AESL_inst_myproject.layer3_out_593_U.if_read & AESL_inst_myproject.layer3_out_593_U.if_empty_n;
    assign fifo_intf_1946.wr_en = AESL_inst_myproject.layer3_out_593_U.if_write & AESL_inst_myproject.layer3_out_593_U.if_full_n;
    assign fifo_intf_1946.fifo_rd_block = 0;
    assign fifo_intf_1946.fifo_wr_block = 0;
    assign fifo_intf_1946.finish = finish;
    csv_file_dump fifo_csv_dumper_1946;
    csv_file_dump cstatus_csv_dumper_1946;
    df_fifo_monitor fifo_monitor_1946;
    df_fifo_intf fifo_intf_1947(clock,reset);
    assign fifo_intf_1947.rd_en = AESL_inst_myproject.layer3_out_594_U.if_read & AESL_inst_myproject.layer3_out_594_U.if_empty_n;
    assign fifo_intf_1947.wr_en = AESL_inst_myproject.layer3_out_594_U.if_write & AESL_inst_myproject.layer3_out_594_U.if_full_n;
    assign fifo_intf_1947.fifo_rd_block = 0;
    assign fifo_intf_1947.fifo_wr_block = 0;
    assign fifo_intf_1947.finish = finish;
    csv_file_dump fifo_csv_dumper_1947;
    csv_file_dump cstatus_csv_dumper_1947;
    df_fifo_monitor fifo_monitor_1947;
    df_fifo_intf fifo_intf_1948(clock,reset);
    assign fifo_intf_1948.rd_en = AESL_inst_myproject.layer3_out_595_U.if_read & AESL_inst_myproject.layer3_out_595_U.if_empty_n;
    assign fifo_intf_1948.wr_en = AESL_inst_myproject.layer3_out_595_U.if_write & AESL_inst_myproject.layer3_out_595_U.if_full_n;
    assign fifo_intf_1948.fifo_rd_block = 0;
    assign fifo_intf_1948.fifo_wr_block = 0;
    assign fifo_intf_1948.finish = finish;
    csv_file_dump fifo_csv_dumper_1948;
    csv_file_dump cstatus_csv_dumper_1948;
    df_fifo_monitor fifo_monitor_1948;
    df_fifo_intf fifo_intf_1949(clock,reset);
    assign fifo_intf_1949.rd_en = AESL_inst_myproject.layer3_out_596_U.if_read & AESL_inst_myproject.layer3_out_596_U.if_empty_n;
    assign fifo_intf_1949.wr_en = AESL_inst_myproject.layer3_out_596_U.if_write & AESL_inst_myproject.layer3_out_596_U.if_full_n;
    assign fifo_intf_1949.fifo_rd_block = 0;
    assign fifo_intf_1949.fifo_wr_block = 0;
    assign fifo_intf_1949.finish = finish;
    csv_file_dump fifo_csv_dumper_1949;
    csv_file_dump cstatus_csv_dumper_1949;
    df_fifo_monitor fifo_monitor_1949;
    df_fifo_intf fifo_intf_1950(clock,reset);
    assign fifo_intf_1950.rd_en = AESL_inst_myproject.layer3_out_597_U.if_read & AESL_inst_myproject.layer3_out_597_U.if_empty_n;
    assign fifo_intf_1950.wr_en = AESL_inst_myproject.layer3_out_597_U.if_write & AESL_inst_myproject.layer3_out_597_U.if_full_n;
    assign fifo_intf_1950.fifo_rd_block = 0;
    assign fifo_intf_1950.fifo_wr_block = 0;
    assign fifo_intf_1950.finish = finish;
    csv_file_dump fifo_csv_dumper_1950;
    csv_file_dump cstatus_csv_dumper_1950;
    df_fifo_monitor fifo_monitor_1950;
    df_fifo_intf fifo_intf_1951(clock,reset);
    assign fifo_intf_1951.rd_en = AESL_inst_myproject.layer3_out_598_U.if_read & AESL_inst_myproject.layer3_out_598_U.if_empty_n;
    assign fifo_intf_1951.wr_en = AESL_inst_myproject.layer3_out_598_U.if_write & AESL_inst_myproject.layer3_out_598_U.if_full_n;
    assign fifo_intf_1951.fifo_rd_block = 0;
    assign fifo_intf_1951.fifo_wr_block = 0;
    assign fifo_intf_1951.finish = finish;
    csv_file_dump fifo_csv_dumper_1951;
    csv_file_dump cstatus_csv_dumper_1951;
    df_fifo_monitor fifo_monitor_1951;
    df_fifo_intf fifo_intf_1952(clock,reset);
    assign fifo_intf_1952.rd_en = AESL_inst_myproject.layer3_out_599_U.if_read & AESL_inst_myproject.layer3_out_599_U.if_empty_n;
    assign fifo_intf_1952.wr_en = AESL_inst_myproject.layer3_out_599_U.if_write & AESL_inst_myproject.layer3_out_599_U.if_full_n;
    assign fifo_intf_1952.fifo_rd_block = 0;
    assign fifo_intf_1952.fifo_wr_block = 0;
    assign fifo_intf_1952.finish = finish;
    csv_file_dump fifo_csv_dumper_1952;
    csv_file_dump cstatus_csv_dumper_1952;
    df_fifo_monitor fifo_monitor_1952;
    df_fifo_intf fifo_intf_1953(clock,reset);
    assign fifo_intf_1953.rd_en = AESL_inst_myproject.layer3_out_600_U.if_read & AESL_inst_myproject.layer3_out_600_U.if_empty_n;
    assign fifo_intf_1953.wr_en = AESL_inst_myproject.layer3_out_600_U.if_write & AESL_inst_myproject.layer3_out_600_U.if_full_n;
    assign fifo_intf_1953.fifo_rd_block = 0;
    assign fifo_intf_1953.fifo_wr_block = 0;
    assign fifo_intf_1953.finish = finish;
    csv_file_dump fifo_csv_dumper_1953;
    csv_file_dump cstatus_csv_dumper_1953;
    df_fifo_monitor fifo_monitor_1953;
    df_fifo_intf fifo_intf_1954(clock,reset);
    assign fifo_intf_1954.rd_en = AESL_inst_myproject.layer3_out_601_U.if_read & AESL_inst_myproject.layer3_out_601_U.if_empty_n;
    assign fifo_intf_1954.wr_en = AESL_inst_myproject.layer3_out_601_U.if_write & AESL_inst_myproject.layer3_out_601_U.if_full_n;
    assign fifo_intf_1954.fifo_rd_block = 0;
    assign fifo_intf_1954.fifo_wr_block = 0;
    assign fifo_intf_1954.finish = finish;
    csv_file_dump fifo_csv_dumper_1954;
    csv_file_dump cstatus_csv_dumper_1954;
    df_fifo_monitor fifo_monitor_1954;
    df_fifo_intf fifo_intf_1955(clock,reset);
    assign fifo_intf_1955.rd_en = AESL_inst_myproject.layer3_out_602_U.if_read & AESL_inst_myproject.layer3_out_602_U.if_empty_n;
    assign fifo_intf_1955.wr_en = AESL_inst_myproject.layer3_out_602_U.if_write & AESL_inst_myproject.layer3_out_602_U.if_full_n;
    assign fifo_intf_1955.fifo_rd_block = 0;
    assign fifo_intf_1955.fifo_wr_block = 0;
    assign fifo_intf_1955.finish = finish;
    csv_file_dump fifo_csv_dumper_1955;
    csv_file_dump cstatus_csv_dumper_1955;
    df_fifo_monitor fifo_monitor_1955;
    df_fifo_intf fifo_intf_1956(clock,reset);
    assign fifo_intf_1956.rd_en = AESL_inst_myproject.layer3_out_603_U.if_read & AESL_inst_myproject.layer3_out_603_U.if_empty_n;
    assign fifo_intf_1956.wr_en = AESL_inst_myproject.layer3_out_603_U.if_write & AESL_inst_myproject.layer3_out_603_U.if_full_n;
    assign fifo_intf_1956.fifo_rd_block = 0;
    assign fifo_intf_1956.fifo_wr_block = 0;
    assign fifo_intf_1956.finish = finish;
    csv_file_dump fifo_csv_dumper_1956;
    csv_file_dump cstatus_csv_dumper_1956;
    df_fifo_monitor fifo_monitor_1956;
    df_fifo_intf fifo_intf_1957(clock,reset);
    assign fifo_intf_1957.rd_en = AESL_inst_myproject.layer3_out_604_U.if_read & AESL_inst_myproject.layer3_out_604_U.if_empty_n;
    assign fifo_intf_1957.wr_en = AESL_inst_myproject.layer3_out_604_U.if_write & AESL_inst_myproject.layer3_out_604_U.if_full_n;
    assign fifo_intf_1957.fifo_rd_block = 0;
    assign fifo_intf_1957.fifo_wr_block = 0;
    assign fifo_intf_1957.finish = finish;
    csv_file_dump fifo_csv_dumper_1957;
    csv_file_dump cstatus_csv_dumper_1957;
    df_fifo_monitor fifo_monitor_1957;
    df_fifo_intf fifo_intf_1958(clock,reset);
    assign fifo_intf_1958.rd_en = AESL_inst_myproject.layer3_out_605_U.if_read & AESL_inst_myproject.layer3_out_605_U.if_empty_n;
    assign fifo_intf_1958.wr_en = AESL_inst_myproject.layer3_out_605_U.if_write & AESL_inst_myproject.layer3_out_605_U.if_full_n;
    assign fifo_intf_1958.fifo_rd_block = 0;
    assign fifo_intf_1958.fifo_wr_block = 0;
    assign fifo_intf_1958.finish = finish;
    csv_file_dump fifo_csv_dumper_1958;
    csv_file_dump cstatus_csv_dumper_1958;
    df_fifo_monitor fifo_monitor_1958;
    df_fifo_intf fifo_intf_1959(clock,reset);
    assign fifo_intf_1959.rd_en = AESL_inst_myproject.layer3_out_606_U.if_read & AESL_inst_myproject.layer3_out_606_U.if_empty_n;
    assign fifo_intf_1959.wr_en = AESL_inst_myproject.layer3_out_606_U.if_write & AESL_inst_myproject.layer3_out_606_U.if_full_n;
    assign fifo_intf_1959.fifo_rd_block = 0;
    assign fifo_intf_1959.fifo_wr_block = 0;
    assign fifo_intf_1959.finish = finish;
    csv_file_dump fifo_csv_dumper_1959;
    csv_file_dump cstatus_csv_dumper_1959;
    df_fifo_monitor fifo_monitor_1959;
    df_fifo_intf fifo_intf_1960(clock,reset);
    assign fifo_intf_1960.rd_en = AESL_inst_myproject.layer3_out_607_U.if_read & AESL_inst_myproject.layer3_out_607_U.if_empty_n;
    assign fifo_intf_1960.wr_en = AESL_inst_myproject.layer3_out_607_U.if_write & AESL_inst_myproject.layer3_out_607_U.if_full_n;
    assign fifo_intf_1960.fifo_rd_block = 0;
    assign fifo_intf_1960.fifo_wr_block = 0;
    assign fifo_intf_1960.finish = finish;
    csv_file_dump fifo_csv_dumper_1960;
    csv_file_dump cstatus_csv_dumper_1960;
    df_fifo_monitor fifo_monitor_1960;
    df_fifo_intf fifo_intf_1961(clock,reset);
    assign fifo_intf_1961.rd_en = AESL_inst_myproject.layer3_out_608_U.if_read & AESL_inst_myproject.layer3_out_608_U.if_empty_n;
    assign fifo_intf_1961.wr_en = AESL_inst_myproject.layer3_out_608_U.if_write & AESL_inst_myproject.layer3_out_608_U.if_full_n;
    assign fifo_intf_1961.fifo_rd_block = 0;
    assign fifo_intf_1961.fifo_wr_block = 0;
    assign fifo_intf_1961.finish = finish;
    csv_file_dump fifo_csv_dumper_1961;
    csv_file_dump cstatus_csv_dumper_1961;
    df_fifo_monitor fifo_monitor_1961;
    df_fifo_intf fifo_intf_1962(clock,reset);
    assign fifo_intf_1962.rd_en = AESL_inst_myproject.layer3_out_609_U.if_read & AESL_inst_myproject.layer3_out_609_U.if_empty_n;
    assign fifo_intf_1962.wr_en = AESL_inst_myproject.layer3_out_609_U.if_write & AESL_inst_myproject.layer3_out_609_U.if_full_n;
    assign fifo_intf_1962.fifo_rd_block = 0;
    assign fifo_intf_1962.fifo_wr_block = 0;
    assign fifo_intf_1962.finish = finish;
    csv_file_dump fifo_csv_dumper_1962;
    csv_file_dump cstatus_csv_dumper_1962;
    df_fifo_monitor fifo_monitor_1962;
    df_fifo_intf fifo_intf_1963(clock,reset);
    assign fifo_intf_1963.rd_en = AESL_inst_myproject.layer3_out_610_U.if_read & AESL_inst_myproject.layer3_out_610_U.if_empty_n;
    assign fifo_intf_1963.wr_en = AESL_inst_myproject.layer3_out_610_U.if_write & AESL_inst_myproject.layer3_out_610_U.if_full_n;
    assign fifo_intf_1963.fifo_rd_block = 0;
    assign fifo_intf_1963.fifo_wr_block = 0;
    assign fifo_intf_1963.finish = finish;
    csv_file_dump fifo_csv_dumper_1963;
    csv_file_dump cstatus_csv_dumper_1963;
    df_fifo_monitor fifo_monitor_1963;
    df_fifo_intf fifo_intf_1964(clock,reset);
    assign fifo_intf_1964.rd_en = AESL_inst_myproject.layer3_out_611_U.if_read & AESL_inst_myproject.layer3_out_611_U.if_empty_n;
    assign fifo_intf_1964.wr_en = AESL_inst_myproject.layer3_out_611_U.if_write & AESL_inst_myproject.layer3_out_611_U.if_full_n;
    assign fifo_intf_1964.fifo_rd_block = 0;
    assign fifo_intf_1964.fifo_wr_block = 0;
    assign fifo_intf_1964.finish = finish;
    csv_file_dump fifo_csv_dumper_1964;
    csv_file_dump cstatus_csv_dumper_1964;
    df_fifo_monitor fifo_monitor_1964;
    df_fifo_intf fifo_intf_1965(clock,reset);
    assign fifo_intf_1965.rd_en = AESL_inst_myproject.layer3_out_612_U.if_read & AESL_inst_myproject.layer3_out_612_U.if_empty_n;
    assign fifo_intf_1965.wr_en = AESL_inst_myproject.layer3_out_612_U.if_write & AESL_inst_myproject.layer3_out_612_U.if_full_n;
    assign fifo_intf_1965.fifo_rd_block = 0;
    assign fifo_intf_1965.fifo_wr_block = 0;
    assign fifo_intf_1965.finish = finish;
    csv_file_dump fifo_csv_dumper_1965;
    csv_file_dump cstatus_csv_dumper_1965;
    df_fifo_monitor fifo_monitor_1965;
    df_fifo_intf fifo_intf_1966(clock,reset);
    assign fifo_intf_1966.rd_en = AESL_inst_myproject.layer3_out_613_U.if_read & AESL_inst_myproject.layer3_out_613_U.if_empty_n;
    assign fifo_intf_1966.wr_en = AESL_inst_myproject.layer3_out_613_U.if_write & AESL_inst_myproject.layer3_out_613_U.if_full_n;
    assign fifo_intf_1966.fifo_rd_block = 0;
    assign fifo_intf_1966.fifo_wr_block = 0;
    assign fifo_intf_1966.finish = finish;
    csv_file_dump fifo_csv_dumper_1966;
    csv_file_dump cstatus_csv_dumper_1966;
    df_fifo_monitor fifo_monitor_1966;
    df_fifo_intf fifo_intf_1967(clock,reset);
    assign fifo_intf_1967.rd_en = AESL_inst_myproject.layer3_out_614_U.if_read & AESL_inst_myproject.layer3_out_614_U.if_empty_n;
    assign fifo_intf_1967.wr_en = AESL_inst_myproject.layer3_out_614_U.if_write & AESL_inst_myproject.layer3_out_614_U.if_full_n;
    assign fifo_intf_1967.fifo_rd_block = 0;
    assign fifo_intf_1967.fifo_wr_block = 0;
    assign fifo_intf_1967.finish = finish;
    csv_file_dump fifo_csv_dumper_1967;
    csv_file_dump cstatus_csv_dumper_1967;
    df_fifo_monitor fifo_monitor_1967;
    df_fifo_intf fifo_intf_1968(clock,reset);
    assign fifo_intf_1968.rd_en = AESL_inst_myproject.layer3_out_615_U.if_read & AESL_inst_myproject.layer3_out_615_U.if_empty_n;
    assign fifo_intf_1968.wr_en = AESL_inst_myproject.layer3_out_615_U.if_write & AESL_inst_myproject.layer3_out_615_U.if_full_n;
    assign fifo_intf_1968.fifo_rd_block = 0;
    assign fifo_intf_1968.fifo_wr_block = 0;
    assign fifo_intf_1968.finish = finish;
    csv_file_dump fifo_csv_dumper_1968;
    csv_file_dump cstatus_csv_dumper_1968;
    df_fifo_monitor fifo_monitor_1968;
    df_fifo_intf fifo_intf_1969(clock,reset);
    assign fifo_intf_1969.rd_en = AESL_inst_myproject.layer3_out_616_U.if_read & AESL_inst_myproject.layer3_out_616_U.if_empty_n;
    assign fifo_intf_1969.wr_en = AESL_inst_myproject.layer3_out_616_U.if_write & AESL_inst_myproject.layer3_out_616_U.if_full_n;
    assign fifo_intf_1969.fifo_rd_block = 0;
    assign fifo_intf_1969.fifo_wr_block = 0;
    assign fifo_intf_1969.finish = finish;
    csv_file_dump fifo_csv_dumper_1969;
    csv_file_dump cstatus_csv_dumper_1969;
    df_fifo_monitor fifo_monitor_1969;
    df_fifo_intf fifo_intf_1970(clock,reset);
    assign fifo_intf_1970.rd_en = AESL_inst_myproject.layer3_out_617_U.if_read & AESL_inst_myproject.layer3_out_617_U.if_empty_n;
    assign fifo_intf_1970.wr_en = AESL_inst_myproject.layer3_out_617_U.if_write & AESL_inst_myproject.layer3_out_617_U.if_full_n;
    assign fifo_intf_1970.fifo_rd_block = 0;
    assign fifo_intf_1970.fifo_wr_block = 0;
    assign fifo_intf_1970.finish = finish;
    csv_file_dump fifo_csv_dumper_1970;
    csv_file_dump cstatus_csv_dumper_1970;
    df_fifo_monitor fifo_monitor_1970;
    df_fifo_intf fifo_intf_1971(clock,reset);
    assign fifo_intf_1971.rd_en = AESL_inst_myproject.layer3_out_618_U.if_read & AESL_inst_myproject.layer3_out_618_U.if_empty_n;
    assign fifo_intf_1971.wr_en = AESL_inst_myproject.layer3_out_618_U.if_write & AESL_inst_myproject.layer3_out_618_U.if_full_n;
    assign fifo_intf_1971.fifo_rd_block = 0;
    assign fifo_intf_1971.fifo_wr_block = 0;
    assign fifo_intf_1971.finish = finish;
    csv_file_dump fifo_csv_dumper_1971;
    csv_file_dump cstatus_csv_dumper_1971;
    df_fifo_monitor fifo_monitor_1971;
    df_fifo_intf fifo_intf_1972(clock,reset);
    assign fifo_intf_1972.rd_en = AESL_inst_myproject.layer3_out_619_U.if_read & AESL_inst_myproject.layer3_out_619_U.if_empty_n;
    assign fifo_intf_1972.wr_en = AESL_inst_myproject.layer3_out_619_U.if_write & AESL_inst_myproject.layer3_out_619_U.if_full_n;
    assign fifo_intf_1972.fifo_rd_block = 0;
    assign fifo_intf_1972.fifo_wr_block = 0;
    assign fifo_intf_1972.finish = finish;
    csv_file_dump fifo_csv_dumper_1972;
    csv_file_dump cstatus_csv_dumper_1972;
    df_fifo_monitor fifo_monitor_1972;
    df_fifo_intf fifo_intf_1973(clock,reset);
    assign fifo_intf_1973.rd_en = AESL_inst_myproject.layer3_out_620_U.if_read & AESL_inst_myproject.layer3_out_620_U.if_empty_n;
    assign fifo_intf_1973.wr_en = AESL_inst_myproject.layer3_out_620_U.if_write & AESL_inst_myproject.layer3_out_620_U.if_full_n;
    assign fifo_intf_1973.fifo_rd_block = 0;
    assign fifo_intf_1973.fifo_wr_block = 0;
    assign fifo_intf_1973.finish = finish;
    csv_file_dump fifo_csv_dumper_1973;
    csv_file_dump cstatus_csv_dumper_1973;
    df_fifo_monitor fifo_monitor_1973;
    df_fifo_intf fifo_intf_1974(clock,reset);
    assign fifo_intf_1974.rd_en = AESL_inst_myproject.layer3_out_621_U.if_read & AESL_inst_myproject.layer3_out_621_U.if_empty_n;
    assign fifo_intf_1974.wr_en = AESL_inst_myproject.layer3_out_621_U.if_write & AESL_inst_myproject.layer3_out_621_U.if_full_n;
    assign fifo_intf_1974.fifo_rd_block = 0;
    assign fifo_intf_1974.fifo_wr_block = 0;
    assign fifo_intf_1974.finish = finish;
    csv_file_dump fifo_csv_dumper_1974;
    csv_file_dump cstatus_csv_dumper_1974;
    df_fifo_monitor fifo_monitor_1974;
    df_fifo_intf fifo_intf_1975(clock,reset);
    assign fifo_intf_1975.rd_en = AESL_inst_myproject.layer3_out_622_U.if_read & AESL_inst_myproject.layer3_out_622_U.if_empty_n;
    assign fifo_intf_1975.wr_en = AESL_inst_myproject.layer3_out_622_U.if_write & AESL_inst_myproject.layer3_out_622_U.if_full_n;
    assign fifo_intf_1975.fifo_rd_block = 0;
    assign fifo_intf_1975.fifo_wr_block = 0;
    assign fifo_intf_1975.finish = finish;
    csv_file_dump fifo_csv_dumper_1975;
    csv_file_dump cstatus_csv_dumper_1975;
    df_fifo_monitor fifo_monitor_1975;
    df_fifo_intf fifo_intf_1976(clock,reset);
    assign fifo_intf_1976.rd_en = AESL_inst_myproject.layer3_out_623_U.if_read & AESL_inst_myproject.layer3_out_623_U.if_empty_n;
    assign fifo_intf_1976.wr_en = AESL_inst_myproject.layer3_out_623_U.if_write & AESL_inst_myproject.layer3_out_623_U.if_full_n;
    assign fifo_intf_1976.fifo_rd_block = 0;
    assign fifo_intf_1976.fifo_wr_block = 0;
    assign fifo_intf_1976.finish = finish;
    csv_file_dump fifo_csv_dumper_1976;
    csv_file_dump cstatus_csv_dumper_1976;
    df_fifo_monitor fifo_monitor_1976;
    df_fifo_intf fifo_intf_1977(clock,reset);
    assign fifo_intf_1977.rd_en = AESL_inst_myproject.layer3_out_624_U.if_read & AESL_inst_myproject.layer3_out_624_U.if_empty_n;
    assign fifo_intf_1977.wr_en = AESL_inst_myproject.layer3_out_624_U.if_write & AESL_inst_myproject.layer3_out_624_U.if_full_n;
    assign fifo_intf_1977.fifo_rd_block = 0;
    assign fifo_intf_1977.fifo_wr_block = 0;
    assign fifo_intf_1977.finish = finish;
    csv_file_dump fifo_csv_dumper_1977;
    csv_file_dump cstatus_csv_dumper_1977;
    df_fifo_monitor fifo_monitor_1977;
    df_fifo_intf fifo_intf_1978(clock,reset);
    assign fifo_intf_1978.rd_en = AESL_inst_myproject.layer3_out_625_U.if_read & AESL_inst_myproject.layer3_out_625_U.if_empty_n;
    assign fifo_intf_1978.wr_en = AESL_inst_myproject.layer3_out_625_U.if_write & AESL_inst_myproject.layer3_out_625_U.if_full_n;
    assign fifo_intf_1978.fifo_rd_block = 0;
    assign fifo_intf_1978.fifo_wr_block = 0;
    assign fifo_intf_1978.finish = finish;
    csv_file_dump fifo_csv_dumper_1978;
    csv_file_dump cstatus_csv_dumper_1978;
    df_fifo_monitor fifo_monitor_1978;
    df_fifo_intf fifo_intf_1979(clock,reset);
    assign fifo_intf_1979.rd_en = AESL_inst_myproject.layer3_out_626_U.if_read & AESL_inst_myproject.layer3_out_626_U.if_empty_n;
    assign fifo_intf_1979.wr_en = AESL_inst_myproject.layer3_out_626_U.if_write & AESL_inst_myproject.layer3_out_626_U.if_full_n;
    assign fifo_intf_1979.fifo_rd_block = 0;
    assign fifo_intf_1979.fifo_wr_block = 0;
    assign fifo_intf_1979.finish = finish;
    csv_file_dump fifo_csv_dumper_1979;
    csv_file_dump cstatus_csv_dumper_1979;
    df_fifo_monitor fifo_monitor_1979;
    df_fifo_intf fifo_intf_1980(clock,reset);
    assign fifo_intf_1980.rd_en = AESL_inst_myproject.layer3_out_627_U.if_read & AESL_inst_myproject.layer3_out_627_U.if_empty_n;
    assign fifo_intf_1980.wr_en = AESL_inst_myproject.layer3_out_627_U.if_write & AESL_inst_myproject.layer3_out_627_U.if_full_n;
    assign fifo_intf_1980.fifo_rd_block = 0;
    assign fifo_intf_1980.fifo_wr_block = 0;
    assign fifo_intf_1980.finish = finish;
    csv_file_dump fifo_csv_dumper_1980;
    csv_file_dump cstatus_csv_dumper_1980;
    df_fifo_monitor fifo_monitor_1980;
    df_fifo_intf fifo_intf_1981(clock,reset);
    assign fifo_intf_1981.rd_en = AESL_inst_myproject.layer3_out_628_U.if_read & AESL_inst_myproject.layer3_out_628_U.if_empty_n;
    assign fifo_intf_1981.wr_en = AESL_inst_myproject.layer3_out_628_U.if_write & AESL_inst_myproject.layer3_out_628_U.if_full_n;
    assign fifo_intf_1981.fifo_rd_block = 0;
    assign fifo_intf_1981.fifo_wr_block = 0;
    assign fifo_intf_1981.finish = finish;
    csv_file_dump fifo_csv_dumper_1981;
    csv_file_dump cstatus_csv_dumper_1981;
    df_fifo_monitor fifo_monitor_1981;
    df_fifo_intf fifo_intf_1982(clock,reset);
    assign fifo_intf_1982.rd_en = AESL_inst_myproject.layer3_out_629_U.if_read & AESL_inst_myproject.layer3_out_629_U.if_empty_n;
    assign fifo_intf_1982.wr_en = AESL_inst_myproject.layer3_out_629_U.if_write & AESL_inst_myproject.layer3_out_629_U.if_full_n;
    assign fifo_intf_1982.fifo_rd_block = 0;
    assign fifo_intf_1982.fifo_wr_block = 0;
    assign fifo_intf_1982.finish = finish;
    csv_file_dump fifo_csv_dumper_1982;
    csv_file_dump cstatus_csv_dumper_1982;
    df_fifo_monitor fifo_monitor_1982;
    df_fifo_intf fifo_intf_1983(clock,reset);
    assign fifo_intf_1983.rd_en = AESL_inst_myproject.layer3_out_630_U.if_read & AESL_inst_myproject.layer3_out_630_U.if_empty_n;
    assign fifo_intf_1983.wr_en = AESL_inst_myproject.layer3_out_630_U.if_write & AESL_inst_myproject.layer3_out_630_U.if_full_n;
    assign fifo_intf_1983.fifo_rd_block = 0;
    assign fifo_intf_1983.fifo_wr_block = 0;
    assign fifo_intf_1983.finish = finish;
    csv_file_dump fifo_csv_dumper_1983;
    csv_file_dump cstatus_csv_dumper_1983;
    df_fifo_monitor fifo_monitor_1983;
    df_fifo_intf fifo_intf_1984(clock,reset);
    assign fifo_intf_1984.rd_en = AESL_inst_myproject.layer3_out_631_U.if_read & AESL_inst_myproject.layer3_out_631_U.if_empty_n;
    assign fifo_intf_1984.wr_en = AESL_inst_myproject.layer3_out_631_U.if_write & AESL_inst_myproject.layer3_out_631_U.if_full_n;
    assign fifo_intf_1984.fifo_rd_block = 0;
    assign fifo_intf_1984.fifo_wr_block = 0;
    assign fifo_intf_1984.finish = finish;
    csv_file_dump fifo_csv_dumper_1984;
    csv_file_dump cstatus_csv_dumper_1984;
    df_fifo_monitor fifo_monitor_1984;
    df_fifo_intf fifo_intf_1985(clock,reset);
    assign fifo_intf_1985.rd_en = AESL_inst_myproject.layer3_out_632_U.if_read & AESL_inst_myproject.layer3_out_632_U.if_empty_n;
    assign fifo_intf_1985.wr_en = AESL_inst_myproject.layer3_out_632_U.if_write & AESL_inst_myproject.layer3_out_632_U.if_full_n;
    assign fifo_intf_1985.fifo_rd_block = 0;
    assign fifo_intf_1985.fifo_wr_block = 0;
    assign fifo_intf_1985.finish = finish;
    csv_file_dump fifo_csv_dumper_1985;
    csv_file_dump cstatus_csv_dumper_1985;
    df_fifo_monitor fifo_monitor_1985;
    df_fifo_intf fifo_intf_1986(clock,reset);
    assign fifo_intf_1986.rd_en = AESL_inst_myproject.layer3_out_633_U.if_read & AESL_inst_myproject.layer3_out_633_U.if_empty_n;
    assign fifo_intf_1986.wr_en = AESL_inst_myproject.layer3_out_633_U.if_write & AESL_inst_myproject.layer3_out_633_U.if_full_n;
    assign fifo_intf_1986.fifo_rd_block = 0;
    assign fifo_intf_1986.fifo_wr_block = 0;
    assign fifo_intf_1986.finish = finish;
    csv_file_dump fifo_csv_dumper_1986;
    csv_file_dump cstatus_csv_dumper_1986;
    df_fifo_monitor fifo_monitor_1986;
    df_fifo_intf fifo_intf_1987(clock,reset);
    assign fifo_intf_1987.rd_en = AESL_inst_myproject.layer3_out_634_U.if_read & AESL_inst_myproject.layer3_out_634_U.if_empty_n;
    assign fifo_intf_1987.wr_en = AESL_inst_myproject.layer3_out_634_U.if_write & AESL_inst_myproject.layer3_out_634_U.if_full_n;
    assign fifo_intf_1987.fifo_rd_block = 0;
    assign fifo_intf_1987.fifo_wr_block = 0;
    assign fifo_intf_1987.finish = finish;
    csv_file_dump fifo_csv_dumper_1987;
    csv_file_dump cstatus_csv_dumper_1987;
    df_fifo_monitor fifo_monitor_1987;
    df_fifo_intf fifo_intf_1988(clock,reset);
    assign fifo_intf_1988.rd_en = AESL_inst_myproject.layer3_out_635_U.if_read & AESL_inst_myproject.layer3_out_635_U.if_empty_n;
    assign fifo_intf_1988.wr_en = AESL_inst_myproject.layer3_out_635_U.if_write & AESL_inst_myproject.layer3_out_635_U.if_full_n;
    assign fifo_intf_1988.fifo_rd_block = 0;
    assign fifo_intf_1988.fifo_wr_block = 0;
    assign fifo_intf_1988.finish = finish;
    csv_file_dump fifo_csv_dumper_1988;
    csv_file_dump cstatus_csv_dumper_1988;
    df_fifo_monitor fifo_monitor_1988;
    df_fifo_intf fifo_intf_1989(clock,reset);
    assign fifo_intf_1989.rd_en = AESL_inst_myproject.layer3_out_636_U.if_read & AESL_inst_myproject.layer3_out_636_U.if_empty_n;
    assign fifo_intf_1989.wr_en = AESL_inst_myproject.layer3_out_636_U.if_write & AESL_inst_myproject.layer3_out_636_U.if_full_n;
    assign fifo_intf_1989.fifo_rd_block = 0;
    assign fifo_intf_1989.fifo_wr_block = 0;
    assign fifo_intf_1989.finish = finish;
    csv_file_dump fifo_csv_dumper_1989;
    csv_file_dump cstatus_csv_dumper_1989;
    df_fifo_monitor fifo_monitor_1989;
    df_fifo_intf fifo_intf_1990(clock,reset);
    assign fifo_intf_1990.rd_en = AESL_inst_myproject.layer3_out_637_U.if_read & AESL_inst_myproject.layer3_out_637_U.if_empty_n;
    assign fifo_intf_1990.wr_en = AESL_inst_myproject.layer3_out_637_U.if_write & AESL_inst_myproject.layer3_out_637_U.if_full_n;
    assign fifo_intf_1990.fifo_rd_block = 0;
    assign fifo_intf_1990.fifo_wr_block = 0;
    assign fifo_intf_1990.finish = finish;
    csv_file_dump fifo_csv_dumper_1990;
    csv_file_dump cstatus_csv_dumper_1990;
    df_fifo_monitor fifo_monitor_1990;
    df_fifo_intf fifo_intf_1991(clock,reset);
    assign fifo_intf_1991.rd_en = AESL_inst_myproject.layer3_out_638_U.if_read & AESL_inst_myproject.layer3_out_638_U.if_empty_n;
    assign fifo_intf_1991.wr_en = AESL_inst_myproject.layer3_out_638_U.if_write & AESL_inst_myproject.layer3_out_638_U.if_full_n;
    assign fifo_intf_1991.fifo_rd_block = 0;
    assign fifo_intf_1991.fifo_wr_block = 0;
    assign fifo_intf_1991.finish = finish;
    csv_file_dump fifo_csv_dumper_1991;
    csv_file_dump cstatus_csv_dumper_1991;
    df_fifo_monitor fifo_monitor_1991;
    df_fifo_intf fifo_intf_1992(clock,reset);
    assign fifo_intf_1992.rd_en = AESL_inst_myproject.layer3_out_639_U.if_read & AESL_inst_myproject.layer3_out_639_U.if_empty_n;
    assign fifo_intf_1992.wr_en = AESL_inst_myproject.layer3_out_639_U.if_write & AESL_inst_myproject.layer3_out_639_U.if_full_n;
    assign fifo_intf_1992.fifo_rd_block = 0;
    assign fifo_intf_1992.fifo_wr_block = 0;
    assign fifo_intf_1992.finish = finish;
    csv_file_dump fifo_csv_dumper_1992;
    csv_file_dump cstatus_csv_dumper_1992;
    df_fifo_monitor fifo_monitor_1992;
    df_fifo_intf fifo_intf_1993(clock,reset);
    assign fifo_intf_1993.rd_en = AESL_inst_myproject.layer3_out_640_U.if_read & AESL_inst_myproject.layer3_out_640_U.if_empty_n;
    assign fifo_intf_1993.wr_en = AESL_inst_myproject.layer3_out_640_U.if_write & AESL_inst_myproject.layer3_out_640_U.if_full_n;
    assign fifo_intf_1993.fifo_rd_block = 0;
    assign fifo_intf_1993.fifo_wr_block = 0;
    assign fifo_intf_1993.finish = finish;
    csv_file_dump fifo_csv_dumper_1993;
    csv_file_dump cstatus_csv_dumper_1993;
    df_fifo_monitor fifo_monitor_1993;
    df_fifo_intf fifo_intf_1994(clock,reset);
    assign fifo_intf_1994.rd_en = AESL_inst_myproject.layer3_out_641_U.if_read & AESL_inst_myproject.layer3_out_641_U.if_empty_n;
    assign fifo_intf_1994.wr_en = AESL_inst_myproject.layer3_out_641_U.if_write & AESL_inst_myproject.layer3_out_641_U.if_full_n;
    assign fifo_intf_1994.fifo_rd_block = 0;
    assign fifo_intf_1994.fifo_wr_block = 0;
    assign fifo_intf_1994.finish = finish;
    csv_file_dump fifo_csv_dumper_1994;
    csv_file_dump cstatus_csv_dumper_1994;
    df_fifo_monitor fifo_monitor_1994;
    df_fifo_intf fifo_intf_1995(clock,reset);
    assign fifo_intf_1995.rd_en = AESL_inst_myproject.layer3_out_642_U.if_read & AESL_inst_myproject.layer3_out_642_U.if_empty_n;
    assign fifo_intf_1995.wr_en = AESL_inst_myproject.layer3_out_642_U.if_write & AESL_inst_myproject.layer3_out_642_U.if_full_n;
    assign fifo_intf_1995.fifo_rd_block = 0;
    assign fifo_intf_1995.fifo_wr_block = 0;
    assign fifo_intf_1995.finish = finish;
    csv_file_dump fifo_csv_dumper_1995;
    csv_file_dump cstatus_csv_dumper_1995;
    df_fifo_monitor fifo_monitor_1995;
    df_fifo_intf fifo_intf_1996(clock,reset);
    assign fifo_intf_1996.rd_en = AESL_inst_myproject.layer3_out_643_U.if_read & AESL_inst_myproject.layer3_out_643_U.if_empty_n;
    assign fifo_intf_1996.wr_en = AESL_inst_myproject.layer3_out_643_U.if_write & AESL_inst_myproject.layer3_out_643_U.if_full_n;
    assign fifo_intf_1996.fifo_rd_block = 0;
    assign fifo_intf_1996.fifo_wr_block = 0;
    assign fifo_intf_1996.finish = finish;
    csv_file_dump fifo_csv_dumper_1996;
    csv_file_dump cstatus_csv_dumper_1996;
    df_fifo_monitor fifo_monitor_1996;
    df_fifo_intf fifo_intf_1997(clock,reset);
    assign fifo_intf_1997.rd_en = AESL_inst_myproject.layer3_out_644_U.if_read & AESL_inst_myproject.layer3_out_644_U.if_empty_n;
    assign fifo_intf_1997.wr_en = AESL_inst_myproject.layer3_out_644_U.if_write & AESL_inst_myproject.layer3_out_644_U.if_full_n;
    assign fifo_intf_1997.fifo_rd_block = 0;
    assign fifo_intf_1997.fifo_wr_block = 0;
    assign fifo_intf_1997.finish = finish;
    csv_file_dump fifo_csv_dumper_1997;
    csv_file_dump cstatus_csv_dumper_1997;
    df_fifo_monitor fifo_monitor_1997;
    df_fifo_intf fifo_intf_1998(clock,reset);
    assign fifo_intf_1998.rd_en = AESL_inst_myproject.layer3_out_645_U.if_read & AESL_inst_myproject.layer3_out_645_U.if_empty_n;
    assign fifo_intf_1998.wr_en = AESL_inst_myproject.layer3_out_645_U.if_write & AESL_inst_myproject.layer3_out_645_U.if_full_n;
    assign fifo_intf_1998.fifo_rd_block = 0;
    assign fifo_intf_1998.fifo_wr_block = 0;
    assign fifo_intf_1998.finish = finish;
    csv_file_dump fifo_csv_dumper_1998;
    csv_file_dump cstatus_csv_dumper_1998;
    df_fifo_monitor fifo_monitor_1998;
    df_fifo_intf fifo_intf_1999(clock,reset);
    assign fifo_intf_1999.rd_en = AESL_inst_myproject.layer3_out_646_U.if_read & AESL_inst_myproject.layer3_out_646_U.if_empty_n;
    assign fifo_intf_1999.wr_en = AESL_inst_myproject.layer3_out_646_U.if_write & AESL_inst_myproject.layer3_out_646_U.if_full_n;
    assign fifo_intf_1999.fifo_rd_block = 0;
    assign fifo_intf_1999.fifo_wr_block = 0;
    assign fifo_intf_1999.finish = finish;
    csv_file_dump fifo_csv_dumper_1999;
    csv_file_dump cstatus_csv_dumper_1999;
    df_fifo_monitor fifo_monitor_1999;
    df_fifo_intf fifo_intf_2000(clock,reset);
    assign fifo_intf_2000.rd_en = AESL_inst_myproject.layer3_out_647_U.if_read & AESL_inst_myproject.layer3_out_647_U.if_empty_n;
    assign fifo_intf_2000.wr_en = AESL_inst_myproject.layer3_out_647_U.if_write & AESL_inst_myproject.layer3_out_647_U.if_full_n;
    assign fifo_intf_2000.fifo_rd_block = 0;
    assign fifo_intf_2000.fifo_wr_block = 0;
    assign fifo_intf_2000.finish = finish;
    csv_file_dump fifo_csv_dumper_2000;
    csv_file_dump cstatus_csv_dumper_2000;
    df_fifo_monitor fifo_monitor_2000;
    df_fifo_intf fifo_intf_2001(clock,reset);
    assign fifo_intf_2001.rd_en = AESL_inst_myproject.layer3_out_648_U.if_read & AESL_inst_myproject.layer3_out_648_U.if_empty_n;
    assign fifo_intf_2001.wr_en = AESL_inst_myproject.layer3_out_648_U.if_write & AESL_inst_myproject.layer3_out_648_U.if_full_n;
    assign fifo_intf_2001.fifo_rd_block = 0;
    assign fifo_intf_2001.fifo_wr_block = 0;
    assign fifo_intf_2001.finish = finish;
    csv_file_dump fifo_csv_dumper_2001;
    csv_file_dump cstatus_csv_dumper_2001;
    df_fifo_monitor fifo_monitor_2001;
    df_fifo_intf fifo_intf_2002(clock,reset);
    assign fifo_intf_2002.rd_en = AESL_inst_myproject.layer3_out_649_U.if_read & AESL_inst_myproject.layer3_out_649_U.if_empty_n;
    assign fifo_intf_2002.wr_en = AESL_inst_myproject.layer3_out_649_U.if_write & AESL_inst_myproject.layer3_out_649_U.if_full_n;
    assign fifo_intf_2002.fifo_rd_block = 0;
    assign fifo_intf_2002.fifo_wr_block = 0;
    assign fifo_intf_2002.finish = finish;
    csv_file_dump fifo_csv_dumper_2002;
    csv_file_dump cstatus_csv_dumper_2002;
    df_fifo_monitor fifo_monitor_2002;
    df_fifo_intf fifo_intf_2003(clock,reset);
    assign fifo_intf_2003.rd_en = AESL_inst_myproject.layer3_out_650_U.if_read & AESL_inst_myproject.layer3_out_650_U.if_empty_n;
    assign fifo_intf_2003.wr_en = AESL_inst_myproject.layer3_out_650_U.if_write & AESL_inst_myproject.layer3_out_650_U.if_full_n;
    assign fifo_intf_2003.fifo_rd_block = 0;
    assign fifo_intf_2003.fifo_wr_block = 0;
    assign fifo_intf_2003.finish = finish;
    csv_file_dump fifo_csv_dumper_2003;
    csv_file_dump cstatus_csv_dumper_2003;
    df_fifo_monitor fifo_monitor_2003;
    df_fifo_intf fifo_intf_2004(clock,reset);
    assign fifo_intf_2004.rd_en = AESL_inst_myproject.layer3_out_651_U.if_read & AESL_inst_myproject.layer3_out_651_U.if_empty_n;
    assign fifo_intf_2004.wr_en = AESL_inst_myproject.layer3_out_651_U.if_write & AESL_inst_myproject.layer3_out_651_U.if_full_n;
    assign fifo_intf_2004.fifo_rd_block = 0;
    assign fifo_intf_2004.fifo_wr_block = 0;
    assign fifo_intf_2004.finish = finish;
    csv_file_dump fifo_csv_dumper_2004;
    csv_file_dump cstatus_csv_dumper_2004;
    df_fifo_monitor fifo_monitor_2004;
    df_fifo_intf fifo_intf_2005(clock,reset);
    assign fifo_intf_2005.rd_en = AESL_inst_myproject.layer3_out_652_U.if_read & AESL_inst_myproject.layer3_out_652_U.if_empty_n;
    assign fifo_intf_2005.wr_en = AESL_inst_myproject.layer3_out_652_U.if_write & AESL_inst_myproject.layer3_out_652_U.if_full_n;
    assign fifo_intf_2005.fifo_rd_block = 0;
    assign fifo_intf_2005.fifo_wr_block = 0;
    assign fifo_intf_2005.finish = finish;
    csv_file_dump fifo_csv_dumper_2005;
    csv_file_dump cstatus_csv_dumper_2005;
    df_fifo_monitor fifo_monitor_2005;
    df_fifo_intf fifo_intf_2006(clock,reset);
    assign fifo_intf_2006.rd_en = AESL_inst_myproject.layer3_out_653_U.if_read & AESL_inst_myproject.layer3_out_653_U.if_empty_n;
    assign fifo_intf_2006.wr_en = AESL_inst_myproject.layer3_out_653_U.if_write & AESL_inst_myproject.layer3_out_653_U.if_full_n;
    assign fifo_intf_2006.fifo_rd_block = 0;
    assign fifo_intf_2006.fifo_wr_block = 0;
    assign fifo_intf_2006.finish = finish;
    csv_file_dump fifo_csv_dumper_2006;
    csv_file_dump cstatus_csv_dumper_2006;
    df_fifo_monitor fifo_monitor_2006;
    df_fifo_intf fifo_intf_2007(clock,reset);
    assign fifo_intf_2007.rd_en = AESL_inst_myproject.layer3_out_654_U.if_read & AESL_inst_myproject.layer3_out_654_U.if_empty_n;
    assign fifo_intf_2007.wr_en = AESL_inst_myproject.layer3_out_654_U.if_write & AESL_inst_myproject.layer3_out_654_U.if_full_n;
    assign fifo_intf_2007.fifo_rd_block = 0;
    assign fifo_intf_2007.fifo_wr_block = 0;
    assign fifo_intf_2007.finish = finish;
    csv_file_dump fifo_csv_dumper_2007;
    csv_file_dump cstatus_csv_dumper_2007;
    df_fifo_monitor fifo_monitor_2007;
    df_fifo_intf fifo_intf_2008(clock,reset);
    assign fifo_intf_2008.rd_en = AESL_inst_myproject.layer3_out_655_U.if_read & AESL_inst_myproject.layer3_out_655_U.if_empty_n;
    assign fifo_intf_2008.wr_en = AESL_inst_myproject.layer3_out_655_U.if_write & AESL_inst_myproject.layer3_out_655_U.if_full_n;
    assign fifo_intf_2008.fifo_rd_block = 0;
    assign fifo_intf_2008.fifo_wr_block = 0;
    assign fifo_intf_2008.finish = finish;
    csv_file_dump fifo_csv_dumper_2008;
    csv_file_dump cstatus_csv_dumper_2008;
    df_fifo_monitor fifo_monitor_2008;
    df_fifo_intf fifo_intf_2009(clock,reset);
    assign fifo_intf_2009.rd_en = AESL_inst_myproject.layer3_out_656_U.if_read & AESL_inst_myproject.layer3_out_656_U.if_empty_n;
    assign fifo_intf_2009.wr_en = AESL_inst_myproject.layer3_out_656_U.if_write & AESL_inst_myproject.layer3_out_656_U.if_full_n;
    assign fifo_intf_2009.fifo_rd_block = 0;
    assign fifo_intf_2009.fifo_wr_block = 0;
    assign fifo_intf_2009.finish = finish;
    csv_file_dump fifo_csv_dumper_2009;
    csv_file_dump cstatus_csv_dumper_2009;
    df_fifo_monitor fifo_monitor_2009;
    df_fifo_intf fifo_intf_2010(clock,reset);
    assign fifo_intf_2010.rd_en = AESL_inst_myproject.layer3_out_657_U.if_read & AESL_inst_myproject.layer3_out_657_U.if_empty_n;
    assign fifo_intf_2010.wr_en = AESL_inst_myproject.layer3_out_657_U.if_write & AESL_inst_myproject.layer3_out_657_U.if_full_n;
    assign fifo_intf_2010.fifo_rd_block = 0;
    assign fifo_intf_2010.fifo_wr_block = 0;
    assign fifo_intf_2010.finish = finish;
    csv_file_dump fifo_csv_dumper_2010;
    csv_file_dump cstatus_csv_dumper_2010;
    df_fifo_monitor fifo_monitor_2010;
    df_fifo_intf fifo_intf_2011(clock,reset);
    assign fifo_intf_2011.rd_en = AESL_inst_myproject.layer3_out_658_U.if_read & AESL_inst_myproject.layer3_out_658_U.if_empty_n;
    assign fifo_intf_2011.wr_en = AESL_inst_myproject.layer3_out_658_U.if_write & AESL_inst_myproject.layer3_out_658_U.if_full_n;
    assign fifo_intf_2011.fifo_rd_block = 0;
    assign fifo_intf_2011.fifo_wr_block = 0;
    assign fifo_intf_2011.finish = finish;
    csv_file_dump fifo_csv_dumper_2011;
    csv_file_dump cstatus_csv_dumper_2011;
    df_fifo_monitor fifo_monitor_2011;
    df_fifo_intf fifo_intf_2012(clock,reset);
    assign fifo_intf_2012.rd_en = AESL_inst_myproject.layer3_out_659_U.if_read & AESL_inst_myproject.layer3_out_659_U.if_empty_n;
    assign fifo_intf_2012.wr_en = AESL_inst_myproject.layer3_out_659_U.if_write & AESL_inst_myproject.layer3_out_659_U.if_full_n;
    assign fifo_intf_2012.fifo_rd_block = 0;
    assign fifo_intf_2012.fifo_wr_block = 0;
    assign fifo_intf_2012.finish = finish;
    csv_file_dump fifo_csv_dumper_2012;
    csv_file_dump cstatus_csv_dumper_2012;
    df_fifo_monitor fifo_monitor_2012;
    df_fifo_intf fifo_intf_2013(clock,reset);
    assign fifo_intf_2013.rd_en = AESL_inst_myproject.layer3_out_660_U.if_read & AESL_inst_myproject.layer3_out_660_U.if_empty_n;
    assign fifo_intf_2013.wr_en = AESL_inst_myproject.layer3_out_660_U.if_write & AESL_inst_myproject.layer3_out_660_U.if_full_n;
    assign fifo_intf_2013.fifo_rd_block = 0;
    assign fifo_intf_2013.fifo_wr_block = 0;
    assign fifo_intf_2013.finish = finish;
    csv_file_dump fifo_csv_dumper_2013;
    csv_file_dump cstatus_csv_dumper_2013;
    df_fifo_monitor fifo_monitor_2013;
    df_fifo_intf fifo_intf_2014(clock,reset);
    assign fifo_intf_2014.rd_en = AESL_inst_myproject.layer3_out_661_U.if_read & AESL_inst_myproject.layer3_out_661_U.if_empty_n;
    assign fifo_intf_2014.wr_en = AESL_inst_myproject.layer3_out_661_U.if_write & AESL_inst_myproject.layer3_out_661_U.if_full_n;
    assign fifo_intf_2014.fifo_rd_block = 0;
    assign fifo_intf_2014.fifo_wr_block = 0;
    assign fifo_intf_2014.finish = finish;
    csv_file_dump fifo_csv_dumper_2014;
    csv_file_dump cstatus_csv_dumper_2014;
    df_fifo_monitor fifo_monitor_2014;
    df_fifo_intf fifo_intf_2015(clock,reset);
    assign fifo_intf_2015.rd_en = AESL_inst_myproject.layer3_out_662_U.if_read & AESL_inst_myproject.layer3_out_662_U.if_empty_n;
    assign fifo_intf_2015.wr_en = AESL_inst_myproject.layer3_out_662_U.if_write & AESL_inst_myproject.layer3_out_662_U.if_full_n;
    assign fifo_intf_2015.fifo_rd_block = 0;
    assign fifo_intf_2015.fifo_wr_block = 0;
    assign fifo_intf_2015.finish = finish;
    csv_file_dump fifo_csv_dumper_2015;
    csv_file_dump cstatus_csv_dumper_2015;
    df_fifo_monitor fifo_monitor_2015;
    df_fifo_intf fifo_intf_2016(clock,reset);
    assign fifo_intf_2016.rd_en = AESL_inst_myproject.layer3_out_663_U.if_read & AESL_inst_myproject.layer3_out_663_U.if_empty_n;
    assign fifo_intf_2016.wr_en = AESL_inst_myproject.layer3_out_663_U.if_write & AESL_inst_myproject.layer3_out_663_U.if_full_n;
    assign fifo_intf_2016.fifo_rd_block = 0;
    assign fifo_intf_2016.fifo_wr_block = 0;
    assign fifo_intf_2016.finish = finish;
    csv_file_dump fifo_csv_dumper_2016;
    csv_file_dump cstatus_csv_dumper_2016;
    df_fifo_monitor fifo_monitor_2016;
    df_fifo_intf fifo_intf_2017(clock,reset);
    assign fifo_intf_2017.rd_en = AESL_inst_myproject.layer3_out_664_U.if_read & AESL_inst_myproject.layer3_out_664_U.if_empty_n;
    assign fifo_intf_2017.wr_en = AESL_inst_myproject.layer3_out_664_U.if_write & AESL_inst_myproject.layer3_out_664_U.if_full_n;
    assign fifo_intf_2017.fifo_rd_block = 0;
    assign fifo_intf_2017.fifo_wr_block = 0;
    assign fifo_intf_2017.finish = finish;
    csv_file_dump fifo_csv_dumper_2017;
    csv_file_dump cstatus_csv_dumper_2017;
    df_fifo_monitor fifo_monitor_2017;
    df_fifo_intf fifo_intf_2018(clock,reset);
    assign fifo_intf_2018.rd_en = AESL_inst_myproject.layer3_out_665_U.if_read & AESL_inst_myproject.layer3_out_665_U.if_empty_n;
    assign fifo_intf_2018.wr_en = AESL_inst_myproject.layer3_out_665_U.if_write & AESL_inst_myproject.layer3_out_665_U.if_full_n;
    assign fifo_intf_2018.fifo_rd_block = 0;
    assign fifo_intf_2018.fifo_wr_block = 0;
    assign fifo_intf_2018.finish = finish;
    csv_file_dump fifo_csv_dumper_2018;
    csv_file_dump cstatus_csv_dumper_2018;
    df_fifo_monitor fifo_monitor_2018;
    df_fifo_intf fifo_intf_2019(clock,reset);
    assign fifo_intf_2019.rd_en = AESL_inst_myproject.layer3_out_666_U.if_read & AESL_inst_myproject.layer3_out_666_U.if_empty_n;
    assign fifo_intf_2019.wr_en = AESL_inst_myproject.layer3_out_666_U.if_write & AESL_inst_myproject.layer3_out_666_U.if_full_n;
    assign fifo_intf_2019.fifo_rd_block = 0;
    assign fifo_intf_2019.fifo_wr_block = 0;
    assign fifo_intf_2019.finish = finish;
    csv_file_dump fifo_csv_dumper_2019;
    csv_file_dump cstatus_csv_dumper_2019;
    df_fifo_monitor fifo_monitor_2019;
    df_fifo_intf fifo_intf_2020(clock,reset);
    assign fifo_intf_2020.rd_en = AESL_inst_myproject.layer3_out_667_U.if_read & AESL_inst_myproject.layer3_out_667_U.if_empty_n;
    assign fifo_intf_2020.wr_en = AESL_inst_myproject.layer3_out_667_U.if_write & AESL_inst_myproject.layer3_out_667_U.if_full_n;
    assign fifo_intf_2020.fifo_rd_block = 0;
    assign fifo_intf_2020.fifo_wr_block = 0;
    assign fifo_intf_2020.finish = finish;
    csv_file_dump fifo_csv_dumper_2020;
    csv_file_dump cstatus_csv_dumper_2020;
    df_fifo_monitor fifo_monitor_2020;
    df_fifo_intf fifo_intf_2021(clock,reset);
    assign fifo_intf_2021.rd_en = AESL_inst_myproject.layer3_out_668_U.if_read & AESL_inst_myproject.layer3_out_668_U.if_empty_n;
    assign fifo_intf_2021.wr_en = AESL_inst_myproject.layer3_out_668_U.if_write & AESL_inst_myproject.layer3_out_668_U.if_full_n;
    assign fifo_intf_2021.fifo_rd_block = 0;
    assign fifo_intf_2021.fifo_wr_block = 0;
    assign fifo_intf_2021.finish = finish;
    csv_file_dump fifo_csv_dumper_2021;
    csv_file_dump cstatus_csv_dumper_2021;
    df_fifo_monitor fifo_monitor_2021;
    df_fifo_intf fifo_intf_2022(clock,reset);
    assign fifo_intf_2022.rd_en = AESL_inst_myproject.layer3_out_669_U.if_read & AESL_inst_myproject.layer3_out_669_U.if_empty_n;
    assign fifo_intf_2022.wr_en = AESL_inst_myproject.layer3_out_669_U.if_write & AESL_inst_myproject.layer3_out_669_U.if_full_n;
    assign fifo_intf_2022.fifo_rd_block = 0;
    assign fifo_intf_2022.fifo_wr_block = 0;
    assign fifo_intf_2022.finish = finish;
    csv_file_dump fifo_csv_dumper_2022;
    csv_file_dump cstatus_csv_dumper_2022;
    df_fifo_monitor fifo_monitor_2022;
    df_fifo_intf fifo_intf_2023(clock,reset);
    assign fifo_intf_2023.rd_en = AESL_inst_myproject.layer3_out_670_U.if_read & AESL_inst_myproject.layer3_out_670_U.if_empty_n;
    assign fifo_intf_2023.wr_en = AESL_inst_myproject.layer3_out_670_U.if_write & AESL_inst_myproject.layer3_out_670_U.if_full_n;
    assign fifo_intf_2023.fifo_rd_block = 0;
    assign fifo_intf_2023.fifo_wr_block = 0;
    assign fifo_intf_2023.finish = finish;
    csv_file_dump fifo_csv_dumper_2023;
    csv_file_dump cstatus_csv_dumper_2023;
    df_fifo_monitor fifo_monitor_2023;
    df_fifo_intf fifo_intf_2024(clock,reset);
    assign fifo_intf_2024.rd_en = AESL_inst_myproject.layer3_out_671_U.if_read & AESL_inst_myproject.layer3_out_671_U.if_empty_n;
    assign fifo_intf_2024.wr_en = AESL_inst_myproject.layer3_out_671_U.if_write & AESL_inst_myproject.layer3_out_671_U.if_full_n;
    assign fifo_intf_2024.fifo_rd_block = 0;
    assign fifo_intf_2024.fifo_wr_block = 0;
    assign fifo_intf_2024.finish = finish;
    csv_file_dump fifo_csv_dumper_2024;
    csv_file_dump cstatus_csv_dumper_2024;
    df_fifo_monitor fifo_monitor_2024;
    df_fifo_intf fifo_intf_2025(clock,reset);
    assign fifo_intf_2025.rd_en = AESL_inst_myproject.layer3_out_672_U.if_read & AESL_inst_myproject.layer3_out_672_U.if_empty_n;
    assign fifo_intf_2025.wr_en = AESL_inst_myproject.layer3_out_672_U.if_write & AESL_inst_myproject.layer3_out_672_U.if_full_n;
    assign fifo_intf_2025.fifo_rd_block = 0;
    assign fifo_intf_2025.fifo_wr_block = 0;
    assign fifo_intf_2025.finish = finish;
    csv_file_dump fifo_csv_dumper_2025;
    csv_file_dump cstatus_csv_dumper_2025;
    df_fifo_monitor fifo_monitor_2025;
    df_fifo_intf fifo_intf_2026(clock,reset);
    assign fifo_intf_2026.rd_en = AESL_inst_myproject.layer3_out_673_U.if_read & AESL_inst_myproject.layer3_out_673_U.if_empty_n;
    assign fifo_intf_2026.wr_en = AESL_inst_myproject.layer3_out_673_U.if_write & AESL_inst_myproject.layer3_out_673_U.if_full_n;
    assign fifo_intf_2026.fifo_rd_block = 0;
    assign fifo_intf_2026.fifo_wr_block = 0;
    assign fifo_intf_2026.finish = finish;
    csv_file_dump fifo_csv_dumper_2026;
    csv_file_dump cstatus_csv_dumper_2026;
    df_fifo_monitor fifo_monitor_2026;
    df_fifo_intf fifo_intf_2027(clock,reset);
    assign fifo_intf_2027.rd_en = AESL_inst_myproject.layer3_out_674_U.if_read & AESL_inst_myproject.layer3_out_674_U.if_empty_n;
    assign fifo_intf_2027.wr_en = AESL_inst_myproject.layer3_out_674_U.if_write & AESL_inst_myproject.layer3_out_674_U.if_full_n;
    assign fifo_intf_2027.fifo_rd_block = 0;
    assign fifo_intf_2027.fifo_wr_block = 0;
    assign fifo_intf_2027.finish = finish;
    csv_file_dump fifo_csv_dumper_2027;
    csv_file_dump cstatus_csv_dumper_2027;
    df_fifo_monitor fifo_monitor_2027;
    df_fifo_intf fifo_intf_2028(clock,reset);
    assign fifo_intf_2028.rd_en = AESL_inst_myproject.layer3_out_675_U.if_read & AESL_inst_myproject.layer3_out_675_U.if_empty_n;
    assign fifo_intf_2028.wr_en = AESL_inst_myproject.layer3_out_675_U.if_write & AESL_inst_myproject.layer3_out_675_U.if_full_n;
    assign fifo_intf_2028.fifo_rd_block = 0;
    assign fifo_intf_2028.fifo_wr_block = 0;
    assign fifo_intf_2028.finish = finish;
    csv_file_dump fifo_csv_dumper_2028;
    csv_file_dump cstatus_csv_dumper_2028;
    df_fifo_monitor fifo_monitor_2028;
    df_fifo_intf fifo_intf_2029(clock,reset);
    assign fifo_intf_2029.rd_en = AESL_inst_myproject.layer3_out_676_U.if_read & AESL_inst_myproject.layer3_out_676_U.if_empty_n;
    assign fifo_intf_2029.wr_en = AESL_inst_myproject.layer3_out_676_U.if_write & AESL_inst_myproject.layer3_out_676_U.if_full_n;
    assign fifo_intf_2029.fifo_rd_block = 0;
    assign fifo_intf_2029.fifo_wr_block = 0;
    assign fifo_intf_2029.finish = finish;
    csv_file_dump fifo_csv_dumper_2029;
    csv_file_dump cstatus_csv_dumper_2029;
    df_fifo_monitor fifo_monitor_2029;
    df_fifo_intf fifo_intf_2030(clock,reset);
    assign fifo_intf_2030.rd_en = AESL_inst_myproject.layer3_out_677_U.if_read & AESL_inst_myproject.layer3_out_677_U.if_empty_n;
    assign fifo_intf_2030.wr_en = AESL_inst_myproject.layer3_out_677_U.if_write & AESL_inst_myproject.layer3_out_677_U.if_full_n;
    assign fifo_intf_2030.fifo_rd_block = 0;
    assign fifo_intf_2030.fifo_wr_block = 0;
    assign fifo_intf_2030.finish = finish;
    csv_file_dump fifo_csv_dumper_2030;
    csv_file_dump cstatus_csv_dumper_2030;
    df_fifo_monitor fifo_monitor_2030;
    df_fifo_intf fifo_intf_2031(clock,reset);
    assign fifo_intf_2031.rd_en = AESL_inst_myproject.layer3_out_678_U.if_read & AESL_inst_myproject.layer3_out_678_U.if_empty_n;
    assign fifo_intf_2031.wr_en = AESL_inst_myproject.layer3_out_678_U.if_write & AESL_inst_myproject.layer3_out_678_U.if_full_n;
    assign fifo_intf_2031.fifo_rd_block = 0;
    assign fifo_intf_2031.fifo_wr_block = 0;
    assign fifo_intf_2031.finish = finish;
    csv_file_dump fifo_csv_dumper_2031;
    csv_file_dump cstatus_csv_dumper_2031;
    df_fifo_monitor fifo_monitor_2031;
    df_fifo_intf fifo_intf_2032(clock,reset);
    assign fifo_intf_2032.rd_en = AESL_inst_myproject.layer3_out_679_U.if_read & AESL_inst_myproject.layer3_out_679_U.if_empty_n;
    assign fifo_intf_2032.wr_en = AESL_inst_myproject.layer3_out_679_U.if_write & AESL_inst_myproject.layer3_out_679_U.if_full_n;
    assign fifo_intf_2032.fifo_rd_block = 0;
    assign fifo_intf_2032.fifo_wr_block = 0;
    assign fifo_intf_2032.finish = finish;
    csv_file_dump fifo_csv_dumper_2032;
    csv_file_dump cstatus_csv_dumper_2032;
    df_fifo_monitor fifo_monitor_2032;
    df_fifo_intf fifo_intf_2033(clock,reset);
    assign fifo_intf_2033.rd_en = AESL_inst_myproject.layer3_out_680_U.if_read & AESL_inst_myproject.layer3_out_680_U.if_empty_n;
    assign fifo_intf_2033.wr_en = AESL_inst_myproject.layer3_out_680_U.if_write & AESL_inst_myproject.layer3_out_680_U.if_full_n;
    assign fifo_intf_2033.fifo_rd_block = 0;
    assign fifo_intf_2033.fifo_wr_block = 0;
    assign fifo_intf_2033.finish = finish;
    csv_file_dump fifo_csv_dumper_2033;
    csv_file_dump cstatus_csv_dumper_2033;
    df_fifo_monitor fifo_monitor_2033;
    df_fifo_intf fifo_intf_2034(clock,reset);
    assign fifo_intf_2034.rd_en = AESL_inst_myproject.layer3_out_681_U.if_read & AESL_inst_myproject.layer3_out_681_U.if_empty_n;
    assign fifo_intf_2034.wr_en = AESL_inst_myproject.layer3_out_681_U.if_write & AESL_inst_myproject.layer3_out_681_U.if_full_n;
    assign fifo_intf_2034.fifo_rd_block = 0;
    assign fifo_intf_2034.fifo_wr_block = 0;
    assign fifo_intf_2034.finish = finish;
    csv_file_dump fifo_csv_dumper_2034;
    csv_file_dump cstatus_csv_dumper_2034;
    df_fifo_monitor fifo_monitor_2034;
    df_fifo_intf fifo_intf_2035(clock,reset);
    assign fifo_intf_2035.rd_en = AESL_inst_myproject.layer3_out_682_U.if_read & AESL_inst_myproject.layer3_out_682_U.if_empty_n;
    assign fifo_intf_2035.wr_en = AESL_inst_myproject.layer3_out_682_U.if_write & AESL_inst_myproject.layer3_out_682_U.if_full_n;
    assign fifo_intf_2035.fifo_rd_block = 0;
    assign fifo_intf_2035.fifo_wr_block = 0;
    assign fifo_intf_2035.finish = finish;
    csv_file_dump fifo_csv_dumper_2035;
    csv_file_dump cstatus_csv_dumper_2035;
    df_fifo_monitor fifo_monitor_2035;
    df_fifo_intf fifo_intf_2036(clock,reset);
    assign fifo_intf_2036.rd_en = AESL_inst_myproject.layer3_out_683_U.if_read & AESL_inst_myproject.layer3_out_683_U.if_empty_n;
    assign fifo_intf_2036.wr_en = AESL_inst_myproject.layer3_out_683_U.if_write & AESL_inst_myproject.layer3_out_683_U.if_full_n;
    assign fifo_intf_2036.fifo_rd_block = 0;
    assign fifo_intf_2036.fifo_wr_block = 0;
    assign fifo_intf_2036.finish = finish;
    csv_file_dump fifo_csv_dumper_2036;
    csv_file_dump cstatus_csv_dumper_2036;
    df_fifo_monitor fifo_monitor_2036;
    df_fifo_intf fifo_intf_2037(clock,reset);
    assign fifo_intf_2037.rd_en = AESL_inst_myproject.layer3_out_684_U.if_read & AESL_inst_myproject.layer3_out_684_U.if_empty_n;
    assign fifo_intf_2037.wr_en = AESL_inst_myproject.layer3_out_684_U.if_write & AESL_inst_myproject.layer3_out_684_U.if_full_n;
    assign fifo_intf_2037.fifo_rd_block = 0;
    assign fifo_intf_2037.fifo_wr_block = 0;
    assign fifo_intf_2037.finish = finish;
    csv_file_dump fifo_csv_dumper_2037;
    csv_file_dump cstatus_csv_dumper_2037;
    df_fifo_monitor fifo_monitor_2037;
    df_fifo_intf fifo_intf_2038(clock,reset);
    assign fifo_intf_2038.rd_en = AESL_inst_myproject.layer3_out_685_U.if_read & AESL_inst_myproject.layer3_out_685_U.if_empty_n;
    assign fifo_intf_2038.wr_en = AESL_inst_myproject.layer3_out_685_U.if_write & AESL_inst_myproject.layer3_out_685_U.if_full_n;
    assign fifo_intf_2038.fifo_rd_block = 0;
    assign fifo_intf_2038.fifo_wr_block = 0;
    assign fifo_intf_2038.finish = finish;
    csv_file_dump fifo_csv_dumper_2038;
    csv_file_dump cstatus_csv_dumper_2038;
    df_fifo_monitor fifo_monitor_2038;
    df_fifo_intf fifo_intf_2039(clock,reset);
    assign fifo_intf_2039.rd_en = AESL_inst_myproject.layer3_out_686_U.if_read & AESL_inst_myproject.layer3_out_686_U.if_empty_n;
    assign fifo_intf_2039.wr_en = AESL_inst_myproject.layer3_out_686_U.if_write & AESL_inst_myproject.layer3_out_686_U.if_full_n;
    assign fifo_intf_2039.fifo_rd_block = 0;
    assign fifo_intf_2039.fifo_wr_block = 0;
    assign fifo_intf_2039.finish = finish;
    csv_file_dump fifo_csv_dumper_2039;
    csv_file_dump cstatus_csv_dumper_2039;
    df_fifo_monitor fifo_monitor_2039;
    df_fifo_intf fifo_intf_2040(clock,reset);
    assign fifo_intf_2040.rd_en = AESL_inst_myproject.layer3_out_687_U.if_read & AESL_inst_myproject.layer3_out_687_U.if_empty_n;
    assign fifo_intf_2040.wr_en = AESL_inst_myproject.layer3_out_687_U.if_write & AESL_inst_myproject.layer3_out_687_U.if_full_n;
    assign fifo_intf_2040.fifo_rd_block = 0;
    assign fifo_intf_2040.fifo_wr_block = 0;
    assign fifo_intf_2040.finish = finish;
    csv_file_dump fifo_csv_dumper_2040;
    csv_file_dump cstatus_csv_dumper_2040;
    df_fifo_monitor fifo_monitor_2040;
    df_fifo_intf fifo_intf_2041(clock,reset);
    assign fifo_intf_2041.rd_en = AESL_inst_myproject.layer3_out_688_U.if_read & AESL_inst_myproject.layer3_out_688_U.if_empty_n;
    assign fifo_intf_2041.wr_en = AESL_inst_myproject.layer3_out_688_U.if_write & AESL_inst_myproject.layer3_out_688_U.if_full_n;
    assign fifo_intf_2041.fifo_rd_block = 0;
    assign fifo_intf_2041.fifo_wr_block = 0;
    assign fifo_intf_2041.finish = finish;
    csv_file_dump fifo_csv_dumper_2041;
    csv_file_dump cstatus_csv_dumper_2041;
    df_fifo_monitor fifo_monitor_2041;
    df_fifo_intf fifo_intf_2042(clock,reset);
    assign fifo_intf_2042.rd_en = AESL_inst_myproject.layer3_out_689_U.if_read & AESL_inst_myproject.layer3_out_689_U.if_empty_n;
    assign fifo_intf_2042.wr_en = AESL_inst_myproject.layer3_out_689_U.if_write & AESL_inst_myproject.layer3_out_689_U.if_full_n;
    assign fifo_intf_2042.fifo_rd_block = 0;
    assign fifo_intf_2042.fifo_wr_block = 0;
    assign fifo_intf_2042.finish = finish;
    csv_file_dump fifo_csv_dumper_2042;
    csv_file_dump cstatus_csv_dumper_2042;
    df_fifo_monitor fifo_monitor_2042;
    df_fifo_intf fifo_intf_2043(clock,reset);
    assign fifo_intf_2043.rd_en = AESL_inst_myproject.layer3_out_690_U.if_read & AESL_inst_myproject.layer3_out_690_U.if_empty_n;
    assign fifo_intf_2043.wr_en = AESL_inst_myproject.layer3_out_690_U.if_write & AESL_inst_myproject.layer3_out_690_U.if_full_n;
    assign fifo_intf_2043.fifo_rd_block = 0;
    assign fifo_intf_2043.fifo_wr_block = 0;
    assign fifo_intf_2043.finish = finish;
    csv_file_dump fifo_csv_dumper_2043;
    csv_file_dump cstatus_csv_dumper_2043;
    df_fifo_monitor fifo_monitor_2043;
    df_fifo_intf fifo_intf_2044(clock,reset);
    assign fifo_intf_2044.rd_en = AESL_inst_myproject.layer3_out_691_U.if_read & AESL_inst_myproject.layer3_out_691_U.if_empty_n;
    assign fifo_intf_2044.wr_en = AESL_inst_myproject.layer3_out_691_U.if_write & AESL_inst_myproject.layer3_out_691_U.if_full_n;
    assign fifo_intf_2044.fifo_rd_block = 0;
    assign fifo_intf_2044.fifo_wr_block = 0;
    assign fifo_intf_2044.finish = finish;
    csv_file_dump fifo_csv_dumper_2044;
    csv_file_dump cstatus_csv_dumper_2044;
    df_fifo_monitor fifo_monitor_2044;
    df_fifo_intf fifo_intf_2045(clock,reset);
    assign fifo_intf_2045.rd_en = AESL_inst_myproject.layer3_out_692_U.if_read & AESL_inst_myproject.layer3_out_692_U.if_empty_n;
    assign fifo_intf_2045.wr_en = AESL_inst_myproject.layer3_out_692_U.if_write & AESL_inst_myproject.layer3_out_692_U.if_full_n;
    assign fifo_intf_2045.fifo_rd_block = 0;
    assign fifo_intf_2045.fifo_wr_block = 0;
    assign fifo_intf_2045.finish = finish;
    csv_file_dump fifo_csv_dumper_2045;
    csv_file_dump cstatus_csv_dumper_2045;
    df_fifo_monitor fifo_monitor_2045;
    df_fifo_intf fifo_intf_2046(clock,reset);
    assign fifo_intf_2046.rd_en = AESL_inst_myproject.layer3_out_693_U.if_read & AESL_inst_myproject.layer3_out_693_U.if_empty_n;
    assign fifo_intf_2046.wr_en = AESL_inst_myproject.layer3_out_693_U.if_write & AESL_inst_myproject.layer3_out_693_U.if_full_n;
    assign fifo_intf_2046.fifo_rd_block = 0;
    assign fifo_intf_2046.fifo_wr_block = 0;
    assign fifo_intf_2046.finish = finish;
    csv_file_dump fifo_csv_dumper_2046;
    csv_file_dump cstatus_csv_dumper_2046;
    df_fifo_monitor fifo_monitor_2046;
    df_fifo_intf fifo_intf_2047(clock,reset);
    assign fifo_intf_2047.rd_en = AESL_inst_myproject.layer3_out_694_U.if_read & AESL_inst_myproject.layer3_out_694_U.if_empty_n;
    assign fifo_intf_2047.wr_en = AESL_inst_myproject.layer3_out_694_U.if_write & AESL_inst_myproject.layer3_out_694_U.if_full_n;
    assign fifo_intf_2047.fifo_rd_block = 0;
    assign fifo_intf_2047.fifo_wr_block = 0;
    assign fifo_intf_2047.finish = finish;
    csv_file_dump fifo_csv_dumper_2047;
    csv_file_dump cstatus_csv_dumper_2047;
    df_fifo_monitor fifo_monitor_2047;
    df_fifo_intf fifo_intf_2048(clock,reset);
    assign fifo_intf_2048.rd_en = AESL_inst_myproject.layer3_out_695_U.if_read & AESL_inst_myproject.layer3_out_695_U.if_empty_n;
    assign fifo_intf_2048.wr_en = AESL_inst_myproject.layer3_out_695_U.if_write & AESL_inst_myproject.layer3_out_695_U.if_full_n;
    assign fifo_intf_2048.fifo_rd_block = 0;
    assign fifo_intf_2048.fifo_wr_block = 0;
    assign fifo_intf_2048.finish = finish;
    csv_file_dump fifo_csv_dumper_2048;
    csv_file_dump cstatus_csv_dumper_2048;
    df_fifo_monitor fifo_monitor_2048;
    df_fifo_intf fifo_intf_2049(clock,reset);
    assign fifo_intf_2049.rd_en = AESL_inst_myproject.layer3_out_696_U.if_read & AESL_inst_myproject.layer3_out_696_U.if_empty_n;
    assign fifo_intf_2049.wr_en = AESL_inst_myproject.layer3_out_696_U.if_write & AESL_inst_myproject.layer3_out_696_U.if_full_n;
    assign fifo_intf_2049.fifo_rd_block = 0;
    assign fifo_intf_2049.fifo_wr_block = 0;
    assign fifo_intf_2049.finish = finish;
    csv_file_dump fifo_csv_dumper_2049;
    csv_file_dump cstatus_csv_dumper_2049;
    df_fifo_monitor fifo_monitor_2049;
    df_fifo_intf fifo_intf_2050(clock,reset);
    assign fifo_intf_2050.rd_en = AESL_inst_myproject.layer3_out_697_U.if_read & AESL_inst_myproject.layer3_out_697_U.if_empty_n;
    assign fifo_intf_2050.wr_en = AESL_inst_myproject.layer3_out_697_U.if_write & AESL_inst_myproject.layer3_out_697_U.if_full_n;
    assign fifo_intf_2050.fifo_rd_block = 0;
    assign fifo_intf_2050.fifo_wr_block = 0;
    assign fifo_intf_2050.finish = finish;
    csv_file_dump fifo_csv_dumper_2050;
    csv_file_dump cstatus_csv_dumper_2050;
    df_fifo_monitor fifo_monitor_2050;
    df_fifo_intf fifo_intf_2051(clock,reset);
    assign fifo_intf_2051.rd_en = AESL_inst_myproject.layer3_out_698_U.if_read & AESL_inst_myproject.layer3_out_698_U.if_empty_n;
    assign fifo_intf_2051.wr_en = AESL_inst_myproject.layer3_out_698_U.if_write & AESL_inst_myproject.layer3_out_698_U.if_full_n;
    assign fifo_intf_2051.fifo_rd_block = 0;
    assign fifo_intf_2051.fifo_wr_block = 0;
    assign fifo_intf_2051.finish = finish;
    csv_file_dump fifo_csv_dumper_2051;
    csv_file_dump cstatus_csv_dumper_2051;
    df_fifo_monitor fifo_monitor_2051;
    df_fifo_intf fifo_intf_2052(clock,reset);
    assign fifo_intf_2052.rd_en = AESL_inst_myproject.layer3_out_699_U.if_read & AESL_inst_myproject.layer3_out_699_U.if_empty_n;
    assign fifo_intf_2052.wr_en = AESL_inst_myproject.layer3_out_699_U.if_write & AESL_inst_myproject.layer3_out_699_U.if_full_n;
    assign fifo_intf_2052.fifo_rd_block = 0;
    assign fifo_intf_2052.fifo_wr_block = 0;
    assign fifo_intf_2052.finish = finish;
    csv_file_dump fifo_csv_dumper_2052;
    csv_file_dump cstatus_csv_dumper_2052;
    df_fifo_monitor fifo_monitor_2052;
    df_fifo_intf fifo_intf_2053(clock,reset);
    assign fifo_intf_2053.rd_en = AESL_inst_myproject.layer3_out_700_U.if_read & AESL_inst_myproject.layer3_out_700_U.if_empty_n;
    assign fifo_intf_2053.wr_en = AESL_inst_myproject.layer3_out_700_U.if_write & AESL_inst_myproject.layer3_out_700_U.if_full_n;
    assign fifo_intf_2053.fifo_rd_block = 0;
    assign fifo_intf_2053.fifo_wr_block = 0;
    assign fifo_intf_2053.finish = finish;
    csv_file_dump fifo_csv_dumper_2053;
    csv_file_dump cstatus_csv_dumper_2053;
    df_fifo_monitor fifo_monitor_2053;
    df_fifo_intf fifo_intf_2054(clock,reset);
    assign fifo_intf_2054.rd_en = AESL_inst_myproject.layer3_out_701_U.if_read & AESL_inst_myproject.layer3_out_701_U.if_empty_n;
    assign fifo_intf_2054.wr_en = AESL_inst_myproject.layer3_out_701_U.if_write & AESL_inst_myproject.layer3_out_701_U.if_full_n;
    assign fifo_intf_2054.fifo_rd_block = 0;
    assign fifo_intf_2054.fifo_wr_block = 0;
    assign fifo_intf_2054.finish = finish;
    csv_file_dump fifo_csv_dumper_2054;
    csv_file_dump cstatus_csv_dumper_2054;
    df_fifo_monitor fifo_monitor_2054;
    df_fifo_intf fifo_intf_2055(clock,reset);
    assign fifo_intf_2055.rd_en = AESL_inst_myproject.layer3_out_702_U.if_read & AESL_inst_myproject.layer3_out_702_U.if_empty_n;
    assign fifo_intf_2055.wr_en = AESL_inst_myproject.layer3_out_702_U.if_write & AESL_inst_myproject.layer3_out_702_U.if_full_n;
    assign fifo_intf_2055.fifo_rd_block = 0;
    assign fifo_intf_2055.fifo_wr_block = 0;
    assign fifo_intf_2055.finish = finish;
    csv_file_dump fifo_csv_dumper_2055;
    csv_file_dump cstatus_csv_dumper_2055;
    df_fifo_monitor fifo_monitor_2055;
    df_fifo_intf fifo_intf_2056(clock,reset);
    assign fifo_intf_2056.rd_en = AESL_inst_myproject.layer3_out_703_U.if_read & AESL_inst_myproject.layer3_out_703_U.if_empty_n;
    assign fifo_intf_2056.wr_en = AESL_inst_myproject.layer3_out_703_U.if_write & AESL_inst_myproject.layer3_out_703_U.if_full_n;
    assign fifo_intf_2056.fifo_rd_block = 0;
    assign fifo_intf_2056.fifo_wr_block = 0;
    assign fifo_intf_2056.finish = finish;
    csv_file_dump fifo_csv_dumper_2056;
    csv_file_dump cstatus_csv_dumper_2056;
    df_fifo_monitor fifo_monitor_2056;
    df_fifo_intf fifo_intf_2057(clock,reset);
    assign fifo_intf_2057.rd_en = AESL_inst_myproject.layer3_out_704_U.if_read & AESL_inst_myproject.layer3_out_704_U.if_empty_n;
    assign fifo_intf_2057.wr_en = AESL_inst_myproject.layer3_out_704_U.if_write & AESL_inst_myproject.layer3_out_704_U.if_full_n;
    assign fifo_intf_2057.fifo_rd_block = 0;
    assign fifo_intf_2057.fifo_wr_block = 0;
    assign fifo_intf_2057.finish = finish;
    csv_file_dump fifo_csv_dumper_2057;
    csv_file_dump cstatus_csv_dumper_2057;
    df_fifo_monitor fifo_monitor_2057;
    df_fifo_intf fifo_intf_2058(clock,reset);
    assign fifo_intf_2058.rd_en = AESL_inst_myproject.layer3_out_705_U.if_read & AESL_inst_myproject.layer3_out_705_U.if_empty_n;
    assign fifo_intf_2058.wr_en = AESL_inst_myproject.layer3_out_705_U.if_write & AESL_inst_myproject.layer3_out_705_U.if_full_n;
    assign fifo_intf_2058.fifo_rd_block = 0;
    assign fifo_intf_2058.fifo_wr_block = 0;
    assign fifo_intf_2058.finish = finish;
    csv_file_dump fifo_csv_dumper_2058;
    csv_file_dump cstatus_csv_dumper_2058;
    df_fifo_monitor fifo_monitor_2058;
    df_fifo_intf fifo_intf_2059(clock,reset);
    assign fifo_intf_2059.rd_en = AESL_inst_myproject.layer3_out_706_U.if_read & AESL_inst_myproject.layer3_out_706_U.if_empty_n;
    assign fifo_intf_2059.wr_en = AESL_inst_myproject.layer3_out_706_U.if_write & AESL_inst_myproject.layer3_out_706_U.if_full_n;
    assign fifo_intf_2059.fifo_rd_block = 0;
    assign fifo_intf_2059.fifo_wr_block = 0;
    assign fifo_intf_2059.finish = finish;
    csv_file_dump fifo_csv_dumper_2059;
    csv_file_dump cstatus_csv_dumper_2059;
    df_fifo_monitor fifo_monitor_2059;
    df_fifo_intf fifo_intf_2060(clock,reset);
    assign fifo_intf_2060.rd_en = AESL_inst_myproject.layer3_out_707_U.if_read & AESL_inst_myproject.layer3_out_707_U.if_empty_n;
    assign fifo_intf_2060.wr_en = AESL_inst_myproject.layer3_out_707_U.if_write & AESL_inst_myproject.layer3_out_707_U.if_full_n;
    assign fifo_intf_2060.fifo_rd_block = 0;
    assign fifo_intf_2060.fifo_wr_block = 0;
    assign fifo_intf_2060.finish = finish;
    csv_file_dump fifo_csv_dumper_2060;
    csv_file_dump cstatus_csv_dumper_2060;
    df_fifo_monitor fifo_monitor_2060;
    df_fifo_intf fifo_intf_2061(clock,reset);
    assign fifo_intf_2061.rd_en = AESL_inst_myproject.layer3_out_708_U.if_read & AESL_inst_myproject.layer3_out_708_U.if_empty_n;
    assign fifo_intf_2061.wr_en = AESL_inst_myproject.layer3_out_708_U.if_write & AESL_inst_myproject.layer3_out_708_U.if_full_n;
    assign fifo_intf_2061.fifo_rd_block = 0;
    assign fifo_intf_2061.fifo_wr_block = 0;
    assign fifo_intf_2061.finish = finish;
    csv_file_dump fifo_csv_dumper_2061;
    csv_file_dump cstatus_csv_dumper_2061;
    df_fifo_monitor fifo_monitor_2061;
    df_fifo_intf fifo_intf_2062(clock,reset);
    assign fifo_intf_2062.rd_en = AESL_inst_myproject.layer3_out_709_U.if_read & AESL_inst_myproject.layer3_out_709_U.if_empty_n;
    assign fifo_intf_2062.wr_en = AESL_inst_myproject.layer3_out_709_U.if_write & AESL_inst_myproject.layer3_out_709_U.if_full_n;
    assign fifo_intf_2062.fifo_rd_block = 0;
    assign fifo_intf_2062.fifo_wr_block = 0;
    assign fifo_intf_2062.finish = finish;
    csv_file_dump fifo_csv_dumper_2062;
    csv_file_dump cstatus_csv_dumper_2062;
    df_fifo_monitor fifo_monitor_2062;
    df_fifo_intf fifo_intf_2063(clock,reset);
    assign fifo_intf_2063.rd_en = AESL_inst_myproject.layer3_out_710_U.if_read & AESL_inst_myproject.layer3_out_710_U.if_empty_n;
    assign fifo_intf_2063.wr_en = AESL_inst_myproject.layer3_out_710_U.if_write & AESL_inst_myproject.layer3_out_710_U.if_full_n;
    assign fifo_intf_2063.fifo_rd_block = 0;
    assign fifo_intf_2063.fifo_wr_block = 0;
    assign fifo_intf_2063.finish = finish;
    csv_file_dump fifo_csv_dumper_2063;
    csv_file_dump cstatus_csv_dumper_2063;
    df_fifo_monitor fifo_monitor_2063;
    df_fifo_intf fifo_intf_2064(clock,reset);
    assign fifo_intf_2064.rd_en = AESL_inst_myproject.layer3_out_711_U.if_read & AESL_inst_myproject.layer3_out_711_U.if_empty_n;
    assign fifo_intf_2064.wr_en = AESL_inst_myproject.layer3_out_711_U.if_write & AESL_inst_myproject.layer3_out_711_U.if_full_n;
    assign fifo_intf_2064.fifo_rd_block = 0;
    assign fifo_intf_2064.fifo_wr_block = 0;
    assign fifo_intf_2064.finish = finish;
    csv_file_dump fifo_csv_dumper_2064;
    csv_file_dump cstatus_csv_dumper_2064;
    df_fifo_monitor fifo_monitor_2064;
    df_fifo_intf fifo_intf_2065(clock,reset);
    assign fifo_intf_2065.rd_en = AESL_inst_myproject.layer3_out_712_U.if_read & AESL_inst_myproject.layer3_out_712_U.if_empty_n;
    assign fifo_intf_2065.wr_en = AESL_inst_myproject.layer3_out_712_U.if_write & AESL_inst_myproject.layer3_out_712_U.if_full_n;
    assign fifo_intf_2065.fifo_rd_block = 0;
    assign fifo_intf_2065.fifo_wr_block = 0;
    assign fifo_intf_2065.finish = finish;
    csv_file_dump fifo_csv_dumper_2065;
    csv_file_dump cstatus_csv_dumper_2065;
    df_fifo_monitor fifo_monitor_2065;
    df_fifo_intf fifo_intf_2066(clock,reset);
    assign fifo_intf_2066.rd_en = AESL_inst_myproject.layer3_out_713_U.if_read & AESL_inst_myproject.layer3_out_713_U.if_empty_n;
    assign fifo_intf_2066.wr_en = AESL_inst_myproject.layer3_out_713_U.if_write & AESL_inst_myproject.layer3_out_713_U.if_full_n;
    assign fifo_intf_2066.fifo_rd_block = 0;
    assign fifo_intf_2066.fifo_wr_block = 0;
    assign fifo_intf_2066.finish = finish;
    csv_file_dump fifo_csv_dumper_2066;
    csv_file_dump cstatus_csv_dumper_2066;
    df_fifo_monitor fifo_monitor_2066;
    df_fifo_intf fifo_intf_2067(clock,reset);
    assign fifo_intf_2067.rd_en = AESL_inst_myproject.layer3_out_714_U.if_read & AESL_inst_myproject.layer3_out_714_U.if_empty_n;
    assign fifo_intf_2067.wr_en = AESL_inst_myproject.layer3_out_714_U.if_write & AESL_inst_myproject.layer3_out_714_U.if_full_n;
    assign fifo_intf_2067.fifo_rd_block = 0;
    assign fifo_intf_2067.fifo_wr_block = 0;
    assign fifo_intf_2067.finish = finish;
    csv_file_dump fifo_csv_dumper_2067;
    csv_file_dump cstatus_csv_dumper_2067;
    df_fifo_monitor fifo_monitor_2067;
    df_fifo_intf fifo_intf_2068(clock,reset);
    assign fifo_intf_2068.rd_en = AESL_inst_myproject.layer3_out_715_U.if_read & AESL_inst_myproject.layer3_out_715_U.if_empty_n;
    assign fifo_intf_2068.wr_en = AESL_inst_myproject.layer3_out_715_U.if_write & AESL_inst_myproject.layer3_out_715_U.if_full_n;
    assign fifo_intf_2068.fifo_rd_block = 0;
    assign fifo_intf_2068.fifo_wr_block = 0;
    assign fifo_intf_2068.finish = finish;
    csv_file_dump fifo_csv_dumper_2068;
    csv_file_dump cstatus_csv_dumper_2068;
    df_fifo_monitor fifo_monitor_2068;
    df_fifo_intf fifo_intf_2069(clock,reset);
    assign fifo_intf_2069.rd_en = AESL_inst_myproject.layer3_out_716_U.if_read & AESL_inst_myproject.layer3_out_716_U.if_empty_n;
    assign fifo_intf_2069.wr_en = AESL_inst_myproject.layer3_out_716_U.if_write & AESL_inst_myproject.layer3_out_716_U.if_full_n;
    assign fifo_intf_2069.fifo_rd_block = 0;
    assign fifo_intf_2069.fifo_wr_block = 0;
    assign fifo_intf_2069.finish = finish;
    csv_file_dump fifo_csv_dumper_2069;
    csv_file_dump cstatus_csv_dumper_2069;
    df_fifo_monitor fifo_monitor_2069;
    df_fifo_intf fifo_intf_2070(clock,reset);
    assign fifo_intf_2070.rd_en = AESL_inst_myproject.layer3_out_717_U.if_read & AESL_inst_myproject.layer3_out_717_U.if_empty_n;
    assign fifo_intf_2070.wr_en = AESL_inst_myproject.layer3_out_717_U.if_write & AESL_inst_myproject.layer3_out_717_U.if_full_n;
    assign fifo_intf_2070.fifo_rd_block = 0;
    assign fifo_intf_2070.fifo_wr_block = 0;
    assign fifo_intf_2070.finish = finish;
    csv_file_dump fifo_csv_dumper_2070;
    csv_file_dump cstatus_csv_dumper_2070;
    df_fifo_monitor fifo_monitor_2070;
    df_fifo_intf fifo_intf_2071(clock,reset);
    assign fifo_intf_2071.rd_en = AESL_inst_myproject.layer3_out_718_U.if_read & AESL_inst_myproject.layer3_out_718_U.if_empty_n;
    assign fifo_intf_2071.wr_en = AESL_inst_myproject.layer3_out_718_U.if_write & AESL_inst_myproject.layer3_out_718_U.if_full_n;
    assign fifo_intf_2071.fifo_rd_block = 0;
    assign fifo_intf_2071.fifo_wr_block = 0;
    assign fifo_intf_2071.finish = finish;
    csv_file_dump fifo_csv_dumper_2071;
    csv_file_dump cstatus_csv_dumper_2071;
    df_fifo_monitor fifo_monitor_2071;
    df_fifo_intf fifo_intf_2072(clock,reset);
    assign fifo_intf_2072.rd_en = AESL_inst_myproject.layer3_out_719_U.if_read & AESL_inst_myproject.layer3_out_719_U.if_empty_n;
    assign fifo_intf_2072.wr_en = AESL_inst_myproject.layer3_out_719_U.if_write & AESL_inst_myproject.layer3_out_719_U.if_full_n;
    assign fifo_intf_2072.fifo_rd_block = 0;
    assign fifo_intf_2072.fifo_wr_block = 0;
    assign fifo_intf_2072.finish = finish;
    csv_file_dump fifo_csv_dumper_2072;
    csv_file_dump cstatus_csv_dumper_2072;
    df_fifo_monitor fifo_monitor_2072;
    df_fifo_intf fifo_intf_2073(clock,reset);
    assign fifo_intf_2073.rd_en = AESL_inst_myproject.layer3_out_720_U.if_read & AESL_inst_myproject.layer3_out_720_U.if_empty_n;
    assign fifo_intf_2073.wr_en = AESL_inst_myproject.layer3_out_720_U.if_write & AESL_inst_myproject.layer3_out_720_U.if_full_n;
    assign fifo_intf_2073.fifo_rd_block = 0;
    assign fifo_intf_2073.fifo_wr_block = 0;
    assign fifo_intf_2073.finish = finish;
    csv_file_dump fifo_csv_dumper_2073;
    csv_file_dump cstatus_csv_dumper_2073;
    df_fifo_monitor fifo_monitor_2073;
    df_fifo_intf fifo_intf_2074(clock,reset);
    assign fifo_intf_2074.rd_en = AESL_inst_myproject.layer3_out_721_U.if_read & AESL_inst_myproject.layer3_out_721_U.if_empty_n;
    assign fifo_intf_2074.wr_en = AESL_inst_myproject.layer3_out_721_U.if_write & AESL_inst_myproject.layer3_out_721_U.if_full_n;
    assign fifo_intf_2074.fifo_rd_block = 0;
    assign fifo_intf_2074.fifo_wr_block = 0;
    assign fifo_intf_2074.finish = finish;
    csv_file_dump fifo_csv_dumper_2074;
    csv_file_dump cstatus_csv_dumper_2074;
    df_fifo_monitor fifo_monitor_2074;
    df_fifo_intf fifo_intf_2075(clock,reset);
    assign fifo_intf_2075.rd_en = AESL_inst_myproject.layer3_out_722_U.if_read & AESL_inst_myproject.layer3_out_722_U.if_empty_n;
    assign fifo_intf_2075.wr_en = AESL_inst_myproject.layer3_out_722_U.if_write & AESL_inst_myproject.layer3_out_722_U.if_full_n;
    assign fifo_intf_2075.fifo_rd_block = 0;
    assign fifo_intf_2075.fifo_wr_block = 0;
    assign fifo_intf_2075.finish = finish;
    csv_file_dump fifo_csv_dumper_2075;
    csv_file_dump cstatus_csv_dumper_2075;
    df_fifo_monitor fifo_monitor_2075;
    df_fifo_intf fifo_intf_2076(clock,reset);
    assign fifo_intf_2076.rd_en = AESL_inst_myproject.layer3_out_723_U.if_read & AESL_inst_myproject.layer3_out_723_U.if_empty_n;
    assign fifo_intf_2076.wr_en = AESL_inst_myproject.layer3_out_723_U.if_write & AESL_inst_myproject.layer3_out_723_U.if_full_n;
    assign fifo_intf_2076.fifo_rd_block = 0;
    assign fifo_intf_2076.fifo_wr_block = 0;
    assign fifo_intf_2076.finish = finish;
    csv_file_dump fifo_csv_dumper_2076;
    csv_file_dump cstatus_csv_dumper_2076;
    df_fifo_monitor fifo_monitor_2076;
    df_fifo_intf fifo_intf_2077(clock,reset);
    assign fifo_intf_2077.rd_en = AESL_inst_myproject.layer3_out_724_U.if_read & AESL_inst_myproject.layer3_out_724_U.if_empty_n;
    assign fifo_intf_2077.wr_en = AESL_inst_myproject.layer3_out_724_U.if_write & AESL_inst_myproject.layer3_out_724_U.if_full_n;
    assign fifo_intf_2077.fifo_rd_block = 0;
    assign fifo_intf_2077.fifo_wr_block = 0;
    assign fifo_intf_2077.finish = finish;
    csv_file_dump fifo_csv_dumper_2077;
    csv_file_dump cstatus_csv_dumper_2077;
    df_fifo_monitor fifo_monitor_2077;
    df_fifo_intf fifo_intf_2078(clock,reset);
    assign fifo_intf_2078.rd_en = AESL_inst_myproject.layer3_out_725_U.if_read & AESL_inst_myproject.layer3_out_725_U.if_empty_n;
    assign fifo_intf_2078.wr_en = AESL_inst_myproject.layer3_out_725_U.if_write & AESL_inst_myproject.layer3_out_725_U.if_full_n;
    assign fifo_intf_2078.fifo_rd_block = 0;
    assign fifo_intf_2078.fifo_wr_block = 0;
    assign fifo_intf_2078.finish = finish;
    csv_file_dump fifo_csv_dumper_2078;
    csv_file_dump cstatus_csv_dumper_2078;
    df_fifo_monitor fifo_monitor_2078;
    df_fifo_intf fifo_intf_2079(clock,reset);
    assign fifo_intf_2079.rd_en = AESL_inst_myproject.layer3_out_726_U.if_read & AESL_inst_myproject.layer3_out_726_U.if_empty_n;
    assign fifo_intf_2079.wr_en = AESL_inst_myproject.layer3_out_726_U.if_write & AESL_inst_myproject.layer3_out_726_U.if_full_n;
    assign fifo_intf_2079.fifo_rd_block = 0;
    assign fifo_intf_2079.fifo_wr_block = 0;
    assign fifo_intf_2079.finish = finish;
    csv_file_dump fifo_csv_dumper_2079;
    csv_file_dump cstatus_csv_dumper_2079;
    df_fifo_monitor fifo_monitor_2079;
    df_fifo_intf fifo_intf_2080(clock,reset);
    assign fifo_intf_2080.rd_en = AESL_inst_myproject.layer3_out_727_U.if_read & AESL_inst_myproject.layer3_out_727_U.if_empty_n;
    assign fifo_intf_2080.wr_en = AESL_inst_myproject.layer3_out_727_U.if_write & AESL_inst_myproject.layer3_out_727_U.if_full_n;
    assign fifo_intf_2080.fifo_rd_block = 0;
    assign fifo_intf_2080.fifo_wr_block = 0;
    assign fifo_intf_2080.finish = finish;
    csv_file_dump fifo_csv_dumper_2080;
    csv_file_dump cstatus_csv_dumper_2080;
    df_fifo_monitor fifo_monitor_2080;
    df_fifo_intf fifo_intf_2081(clock,reset);
    assign fifo_intf_2081.rd_en = AESL_inst_myproject.layer3_out_728_U.if_read & AESL_inst_myproject.layer3_out_728_U.if_empty_n;
    assign fifo_intf_2081.wr_en = AESL_inst_myproject.layer3_out_728_U.if_write & AESL_inst_myproject.layer3_out_728_U.if_full_n;
    assign fifo_intf_2081.fifo_rd_block = 0;
    assign fifo_intf_2081.fifo_wr_block = 0;
    assign fifo_intf_2081.finish = finish;
    csv_file_dump fifo_csv_dumper_2081;
    csv_file_dump cstatus_csv_dumper_2081;
    df_fifo_monitor fifo_monitor_2081;
    df_fifo_intf fifo_intf_2082(clock,reset);
    assign fifo_intf_2082.rd_en = AESL_inst_myproject.layer3_out_729_U.if_read & AESL_inst_myproject.layer3_out_729_U.if_empty_n;
    assign fifo_intf_2082.wr_en = AESL_inst_myproject.layer3_out_729_U.if_write & AESL_inst_myproject.layer3_out_729_U.if_full_n;
    assign fifo_intf_2082.fifo_rd_block = 0;
    assign fifo_intf_2082.fifo_wr_block = 0;
    assign fifo_intf_2082.finish = finish;
    csv_file_dump fifo_csv_dumper_2082;
    csv_file_dump cstatus_csv_dumper_2082;
    df_fifo_monitor fifo_monitor_2082;
    df_fifo_intf fifo_intf_2083(clock,reset);
    assign fifo_intf_2083.rd_en = AESL_inst_myproject.layer3_out_730_U.if_read & AESL_inst_myproject.layer3_out_730_U.if_empty_n;
    assign fifo_intf_2083.wr_en = AESL_inst_myproject.layer3_out_730_U.if_write & AESL_inst_myproject.layer3_out_730_U.if_full_n;
    assign fifo_intf_2083.fifo_rd_block = 0;
    assign fifo_intf_2083.fifo_wr_block = 0;
    assign fifo_intf_2083.finish = finish;
    csv_file_dump fifo_csv_dumper_2083;
    csv_file_dump cstatus_csv_dumper_2083;
    df_fifo_monitor fifo_monitor_2083;
    df_fifo_intf fifo_intf_2084(clock,reset);
    assign fifo_intf_2084.rd_en = AESL_inst_myproject.layer3_out_731_U.if_read & AESL_inst_myproject.layer3_out_731_U.if_empty_n;
    assign fifo_intf_2084.wr_en = AESL_inst_myproject.layer3_out_731_U.if_write & AESL_inst_myproject.layer3_out_731_U.if_full_n;
    assign fifo_intf_2084.fifo_rd_block = 0;
    assign fifo_intf_2084.fifo_wr_block = 0;
    assign fifo_intf_2084.finish = finish;
    csv_file_dump fifo_csv_dumper_2084;
    csv_file_dump cstatus_csv_dumper_2084;
    df_fifo_monitor fifo_monitor_2084;
    df_fifo_intf fifo_intf_2085(clock,reset);
    assign fifo_intf_2085.rd_en = AESL_inst_myproject.layer3_out_732_U.if_read & AESL_inst_myproject.layer3_out_732_U.if_empty_n;
    assign fifo_intf_2085.wr_en = AESL_inst_myproject.layer3_out_732_U.if_write & AESL_inst_myproject.layer3_out_732_U.if_full_n;
    assign fifo_intf_2085.fifo_rd_block = 0;
    assign fifo_intf_2085.fifo_wr_block = 0;
    assign fifo_intf_2085.finish = finish;
    csv_file_dump fifo_csv_dumper_2085;
    csv_file_dump cstatus_csv_dumper_2085;
    df_fifo_monitor fifo_monitor_2085;
    df_fifo_intf fifo_intf_2086(clock,reset);
    assign fifo_intf_2086.rd_en = AESL_inst_myproject.layer3_out_733_U.if_read & AESL_inst_myproject.layer3_out_733_U.if_empty_n;
    assign fifo_intf_2086.wr_en = AESL_inst_myproject.layer3_out_733_U.if_write & AESL_inst_myproject.layer3_out_733_U.if_full_n;
    assign fifo_intf_2086.fifo_rd_block = 0;
    assign fifo_intf_2086.fifo_wr_block = 0;
    assign fifo_intf_2086.finish = finish;
    csv_file_dump fifo_csv_dumper_2086;
    csv_file_dump cstatus_csv_dumper_2086;
    df_fifo_monitor fifo_monitor_2086;
    df_fifo_intf fifo_intf_2087(clock,reset);
    assign fifo_intf_2087.rd_en = AESL_inst_myproject.layer3_out_734_U.if_read & AESL_inst_myproject.layer3_out_734_U.if_empty_n;
    assign fifo_intf_2087.wr_en = AESL_inst_myproject.layer3_out_734_U.if_write & AESL_inst_myproject.layer3_out_734_U.if_full_n;
    assign fifo_intf_2087.fifo_rd_block = 0;
    assign fifo_intf_2087.fifo_wr_block = 0;
    assign fifo_intf_2087.finish = finish;
    csv_file_dump fifo_csv_dumper_2087;
    csv_file_dump cstatus_csv_dumper_2087;
    df_fifo_monitor fifo_monitor_2087;
    df_fifo_intf fifo_intf_2088(clock,reset);
    assign fifo_intf_2088.rd_en = AESL_inst_myproject.layer3_out_735_U.if_read & AESL_inst_myproject.layer3_out_735_U.if_empty_n;
    assign fifo_intf_2088.wr_en = AESL_inst_myproject.layer3_out_735_U.if_write & AESL_inst_myproject.layer3_out_735_U.if_full_n;
    assign fifo_intf_2088.fifo_rd_block = 0;
    assign fifo_intf_2088.fifo_wr_block = 0;
    assign fifo_intf_2088.finish = finish;
    csv_file_dump fifo_csv_dumper_2088;
    csv_file_dump cstatus_csv_dumper_2088;
    df_fifo_monitor fifo_monitor_2088;
    df_fifo_intf fifo_intf_2089(clock,reset);
    assign fifo_intf_2089.rd_en = AESL_inst_myproject.layer3_out_736_U.if_read & AESL_inst_myproject.layer3_out_736_U.if_empty_n;
    assign fifo_intf_2089.wr_en = AESL_inst_myproject.layer3_out_736_U.if_write & AESL_inst_myproject.layer3_out_736_U.if_full_n;
    assign fifo_intf_2089.fifo_rd_block = 0;
    assign fifo_intf_2089.fifo_wr_block = 0;
    assign fifo_intf_2089.finish = finish;
    csv_file_dump fifo_csv_dumper_2089;
    csv_file_dump cstatus_csv_dumper_2089;
    df_fifo_monitor fifo_monitor_2089;
    df_fifo_intf fifo_intf_2090(clock,reset);
    assign fifo_intf_2090.rd_en = AESL_inst_myproject.layer3_out_737_U.if_read & AESL_inst_myproject.layer3_out_737_U.if_empty_n;
    assign fifo_intf_2090.wr_en = AESL_inst_myproject.layer3_out_737_U.if_write & AESL_inst_myproject.layer3_out_737_U.if_full_n;
    assign fifo_intf_2090.fifo_rd_block = 0;
    assign fifo_intf_2090.fifo_wr_block = 0;
    assign fifo_intf_2090.finish = finish;
    csv_file_dump fifo_csv_dumper_2090;
    csv_file_dump cstatus_csv_dumper_2090;
    df_fifo_monitor fifo_monitor_2090;
    df_fifo_intf fifo_intf_2091(clock,reset);
    assign fifo_intf_2091.rd_en = AESL_inst_myproject.layer3_out_738_U.if_read & AESL_inst_myproject.layer3_out_738_U.if_empty_n;
    assign fifo_intf_2091.wr_en = AESL_inst_myproject.layer3_out_738_U.if_write & AESL_inst_myproject.layer3_out_738_U.if_full_n;
    assign fifo_intf_2091.fifo_rd_block = 0;
    assign fifo_intf_2091.fifo_wr_block = 0;
    assign fifo_intf_2091.finish = finish;
    csv_file_dump fifo_csv_dumper_2091;
    csv_file_dump cstatus_csv_dumper_2091;
    df_fifo_monitor fifo_monitor_2091;
    df_fifo_intf fifo_intf_2092(clock,reset);
    assign fifo_intf_2092.rd_en = AESL_inst_myproject.layer3_out_739_U.if_read & AESL_inst_myproject.layer3_out_739_U.if_empty_n;
    assign fifo_intf_2092.wr_en = AESL_inst_myproject.layer3_out_739_U.if_write & AESL_inst_myproject.layer3_out_739_U.if_full_n;
    assign fifo_intf_2092.fifo_rd_block = 0;
    assign fifo_intf_2092.fifo_wr_block = 0;
    assign fifo_intf_2092.finish = finish;
    csv_file_dump fifo_csv_dumper_2092;
    csv_file_dump cstatus_csv_dumper_2092;
    df_fifo_monitor fifo_monitor_2092;
    df_fifo_intf fifo_intf_2093(clock,reset);
    assign fifo_intf_2093.rd_en = AESL_inst_myproject.layer3_out_740_U.if_read & AESL_inst_myproject.layer3_out_740_U.if_empty_n;
    assign fifo_intf_2093.wr_en = AESL_inst_myproject.layer3_out_740_U.if_write & AESL_inst_myproject.layer3_out_740_U.if_full_n;
    assign fifo_intf_2093.fifo_rd_block = 0;
    assign fifo_intf_2093.fifo_wr_block = 0;
    assign fifo_intf_2093.finish = finish;
    csv_file_dump fifo_csv_dumper_2093;
    csv_file_dump cstatus_csv_dumper_2093;
    df_fifo_monitor fifo_monitor_2093;
    df_fifo_intf fifo_intf_2094(clock,reset);
    assign fifo_intf_2094.rd_en = AESL_inst_myproject.layer3_out_741_U.if_read & AESL_inst_myproject.layer3_out_741_U.if_empty_n;
    assign fifo_intf_2094.wr_en = AESL_inst_myproject.layer3_out_741_U.if_write & AESL_inst_myproject.layer3_out_741_U.if_full_n;
    assign fifo_intf_2094.fifo_rd_block = 0;
    assign fifo_intf_2094.fifo_wr_block = 0;
    assign fifo_intf_2094.finish = finish;
    csv_file_dump fifo_csv_dumper_2094;
    csv_file_dump cstatus_csv_dumper_2094;
    df_fifo_monitor fifo_monitor_2094;
    df_fifo_intf fifo_intf_2095(clock,reset);
    assign fifo_intf_2095.rd_en = AESL_inst_myproject.layer3_out_742_U.if_read & AESL_inst_myproject.layer3_out_742_U.if_empty_n;
    assign fifo_intf_2095.wr_en = AESL_inst_myproject.layer3_out_742_U.if_write & AESL_inst_myproject.layer3_out_742_U.if_full_n;
    assign fifo_intf_2095.fifo_rd_block = 0;
    assign fifo_intf_2095.fifo_wr_block = 0;
    assign fifo_intf_2095.finish = finish;
    csv_file_dump fifo_csv_dumper_2095;
    csv_file_dump cstatus_csv_dumper_2095;
    df_fifo_monitor fifo_monitor_2095;
    df_fifo_intf fifo_intf_2096(clock,reset);
    assign fifo_intf_2096.rd_en = AESL_inst_myproject.layer3_out_743_U.if_read & AESL_inst_myproject.layer3_out_743_U.if_empty_n;
    assign fifo_intf_2096.wr_en = AESL_inst_myproject.layer3_out_743_U.if_write & AESL_inst_myproject.layer3_out_743_U.if_full_n;
    assign fifo_intf_2096.fifo_rd_block = 0;
    assign fifo_intf_2096.fifo_wr_block = 0;
    assign fifo_intf_2096.finish = finish;
    csv_file_dump fifo_csv_dumper_2096;
    csv_file_dump cstatus_csv_dumper_2096;
    df_fifo_monitor fifo_monitor_2096;
    df_fifo_intf fifo_intf_2097(clock,reset);
    assign fifo_intf_2097.rd_en = AESL_inst_myproject.layer3_out_744_U.if_read & AESL_inst_myproject.layer3_out_744_U.if_empty_n;
    assign fifo_intf_2097.wr_en = AESL_inst_myproject.layer3_out_744_U.if_write & AESL_inst_myproject.layer3_out_744_U.if_full_n;
    assign fifo_intf_2097.fifo_rd_block = 0;
    assign fifo_intf_2097.fifo_wr_block = 0;
    assign fifo_intf_2097.finish = finish;
    csv_file_dump fifo_csv_dumper_2097;
    csv_file_dump cstatus_csv_dumper_2097;
    df_fifo_monitor fifo_monitor_2097;
    df_fifo_intf fifo_intf_2098(clock,reset);
    assign fifo_intf_2098.rd_en = AESL_inst_myproject.layer3_out_745_U.if_read & AESL_inst_myproject.layer3_out_745_U.if_empty_n;
    assign fifo_intf_2098.wr_en = AESL_inst_myproject.layer3_out_745_U.if_write & AESL_inst_myproject.layer3_out_745_U.if_full_n;
    assign fifo_intf_2098.fifo_rd_block = 0;
    assign fifo_intf_2098.fifo_wr_block = 0;
    assign fifo_intf_2098.finish = finish;
    csv_file_dump fifo_csv_dumper_2098;
    csv_file_dump cstatus_csv_dumper_2098;
    df_fifo_monitor fifo_monitor_2098;
    df_fifo_intf fifo_intf_2099(clock,reset);
    assign fifo_intf_2099.rd_en = AESL_inst_myproject.layer3_out_746_U.if_read & AESL_inst_myproject.layer3_out_746_U.if_empty_n;
    assign fifo_intf_2099.wr_en = AESL_inst_myproject.layer3_out_746_U.if_write & AESL_inst_myproject.layer3_out_746_U.if_full_n;
    assign fifo_intf_2099.fifo_rd_block = 0;
    assign fifo_intf_2099.fifo_wr_block = 0;
    assign fifo_intf_2099.finish = finish;
    csv_file_dump fifo_csv_dumper_2099;
    csv_file_dump cstatus_csv_dumper_2099;
    df_fifo_monitor fifo_monitor_2099;
    df_fifo_intf fifo_intf_2100(clock,reset);
    assign fifo_intf_2100.rd_en = AESL_inst_myproject.layer3_out_747_U.if_read & AESL_inst_myproject.layer3_out_747_U.if_empty_n;
    assign fifo_intf_2100.wr_en = AESL_inst_myproject.layer3_out_747_U.if_write & AESL_inst_myproject.layer3_out_747_U.if_full_n;
    assign fifo_intf_2100.fifo_rd_block = 0;
    assign fifo_intf_2100.fifo_wr_block = 0;
    assign fifo_intf_2100.finish = finish;
    csv_file_dump fifo_csv_dumper_2100;
    csv_file_dump cstatus_csv_dumper_2100;
    df_fifo_monitor fifo_monitor_2100;
    df_fifo_intf fifo_intf_2101(clock,reset);
    assign fifo_intf_2101.rd_en = AESL_inst_myproject.layer3_out_748_U.if_read & AESL_inst_myproject.layer3_out_748_U.if_empty_n;
    assign fifo_intf_2101.wr_en = AESL_inst_myproject.layer3_out_748_U.if_write & AESL_inst_myproject.layer3_out_748_U.if_full_n;
    assign fifo_intf_2101.fifo_rd_block = 0;
    assign fifo_intf_2101.fifo_wr_block = 0;
    assign fifo_intf_2101.finish = finish;
    csv_file_dump fifo_csv_dumper_2101;
    csv_file_dump cstatus_csv_dumper_2101;
    df_fifo_monitor fifo_monitor_2101;
    df_fifo_intf fifo_intf_2102(clock,reset);
    assign fifo_intf_2102.rd_en = AESL_inst_myproject.layer3_out_749_U.if_read & AESL_inst_myproject.layer3_out_749_U.if_empty_n;
    assign fifo_intf_2102.wr_en = AESL_inst_myproject.layer3_out_749_U.if_write & AESL_inst_myproject.layer3_out_749_U.if_full_n;
    assign fifo_intf_2102.fifo_rd_block = 0;
    assign fifo_intf_2102.fifo_wr_block = 0;
    assign fifo_intf_2102.finish = finish;
    csv_file_dump fifo_csv_dumper_2102;
    csv_file_dump cstatus_csv_dumper_2102;
    df_fifo_monitor fifo_monitor_2102;
    df_fifo_intf fifo_intf_2103(clock,reset);
    assign fifo_intf_2103.rd_en = AESL_inst_myproject.layer3_out_750_U.if_read & AESL_inst_myproject.layer3_out_750_U.if_empty_n;
    assign fifo_intf_2103.wr_en = AESL_inst_myproject.layer3_out_750_U.if_write & AESL_inst_myproject.layer3_out_750_U.if_full_n;
    assign fifo_intf_2103.fifo_rd_block = 0;
    assign fifo_intf_2103.fifo_wr_block = 0;
    assign fifo_intf_2103.finish = finish;
    csv_file_dump fifo_csv_dumper_2103;
    csv_file_dump cstatus_csv_dumper_2103;
    df_fifo_monitor fifo_monitor_2103;
    df_fifo_intf fifo_intf_2104(clock,reset);
    assign fifo_intf_2104.rd_en = AESL_inst_myproject.layer3_out_751_U.if_read & AESL_inst_myproject.layer3_out_751_U.if_empty_n;
    assign fifo_intf_2104.wr_en = AESL_inst_myproject.layer3_out_751_U.if_write & AESL_inst_myproject.layer3_out_751_U.if_full_n;
    assign fifo_intf_2104.fifo_rd_block = 0;
    assign fifo_intf_2104.fifo_wr_block = 0;
    assign fifo_intf_2104.finish = finish;
    csv_file_dump fifo_csv_dumper_2104;
    csv_file_dump cstatus_csv_dumper_2104;
    df_fifo_monitor fifo_monitor_2104;
    df_fifo_intf fifo_intf_2105(clock,reset);
    assign fifo_intf_2105.rd_en = AESL_inst_myproject.layer3_out_752_U.if_read & AESL_inst_myproject.layer3_out_752_U.if_empty_n;
    assign fifo_intf_2105.wr_en = AESL_inst_myproject.layer3_out_752_U.if_write & AESL_inst_myproject.layer3_out_752_U.if_full_n;
    assign fifo_intf_2105.fifo_rd_block = 0;
    assign fifo_intf_2105.fifo_wr_block = 0;
    assign fifo_intf_2105.finish = finish;
    csv_file_dump fifo_csv_dumper_2105;
    csv_file_dump cstatus_csv_dumper_2105;
    df_fifo_monitor fifo_monitor_2105;
    df_fifo_intf fifo_intf_2106(clock,reset);
    assign fifo_intf_2106.rd_en = AESL_inst_myproject.layer3_out_753_U.if_read & AESL_inst_myproject.layer3_out_753_U.if_empty_n;
    assign fifo_intf_2106.wr_en = AESL_inst_myproject.layer3_out_753_U.if_write & AESL_inst_myproject.layer3_out_753_U.if_full_n;
    assign fifo_intf_2106.fifo_rd_block = 0;
    assign fifo_intf_2106.fifo_wr_block = 0;
    assign fifo_intf_2106.finish = finish;
    csv_file_dump fifo_csv_dumper_2106;
    csv_file_dump cstatus_csv_dumper_2106;
    df_fifo_monitor fifo_monitor_2106;
    df_fifo_intf fifo_intf_2107(clock,reset);
    assign fifo_intf_2107.rd_en = AESL_inst_myproject.layer3_out_754_U.if_read & AESL_inst_myproject.layer3_out_754_U.if_empty_n;
    assign fifo_intf_2107.wr_en = AESL_inst_myproject.layer3_out_754_U.if_write & AESL_inst_myproject.layer3_out_754_U.if_full_n;
    assign fifo_intf_2107.fifo_rd_block = 0;
    assign fifo_intf_2107.fifo_wr_block = 0;
    assign fifo_intf_2107.finish = finish;
    csv_file_dump fifo_csv_dumper_2107;
    csv_file_dump cstatus_csv_dumper_2107;
    df_fifo_monitor fifo_monitor_2107;
    df_fifo_intf fifo_intf_2108(clock,reset);
    assign fifo_intf_2108.rd_en = AESL_inst_myproject.layer3_out_755_U.if_read & AESL_inst_myproject.layer3_out_755_U.if_empty_n;
    assign fifo_intf_2108.wr_en = AESL_inst_myproject.layer3_out_755_U.if_write & AESL_inst_myproject.layer3_out_755_U.if_full_n;
    assign fifo_intf_2108.fifo_rd_block = 0;
    assign fifo_intf_2108.fifo_wr_block = 0;
    assign fifo_intf_2108.finish = finish;
    csv_file_dump fifo_csv_dumper_2108;
    csv_file_dump cstatus_csv_dumper_2108;
    df_fifo_monitor fifo_monitor_2108;
    df_fifo_intf fifo_intf_2109(clock,reset);
    assign fifo_intf_2109.rd_en = AESL_inst_myproject.layer3_out_756_U.if_read & AESL_inst_myproject.layer3_out_756_U.if_empty_n;
    assign fifo_intf_2109.wr_en = AESL_inst_myproject.layer3_out_756_U.if_write & AESL_inst_myproject.layer3_out_756_U.if_full_n;
    assign fifo_intf_2109.fifo_rd_block = 0;
    assign fifo_intf_2109.fifo_wr_block = 0;
    assign fifo_intf_2109.finish = finish;
    csv_file_dump fifo_csv_dumper_2109;
    csv_file_dump cstatus_csv_dumper_2109;
    df_fifo_monitor fifo_monitor_2109;
    df_fifo_intf fifo_intf_2110(clock,reset);
    assign fifo_intf_2110.rd_en = AESL_inst_myproject.layer3_out_757_U.if_read & AESL_inst_myproject.layer3_out_757_U.if_empty_n;
    assign fifo_intf_2110.wr_en = AESL_inst_myproject.layer3_out_757_U.if_write & AESL_inst_myproject.layer3_out_757_U.if_full_n;
    assign fifo_intf_2110.fifo_rd_block = 0;
    assign fifo_intf_2110.fifo_wr_block = 0;
    assign fifo_intf_2110.finish = finish;
    csv_file_dump fifo_csv_dumper_2110;
    csv_file_dump cstatus_csv_dumper_2110;
    df_fifo_monitor fifo_monitor_2110;
    df_fifo_intf fifo_intf_2111(clock,reset);
    assign fifo_intf_2111.rd_en = AESL_inst_myproject.layer3_out_758_U.if_read & AESL_inst_myproject.layer3_out_758_U.if_empty_n;
    assign fifo_intf_2111.wr_en = AESL_inst_myproject.layer3_out_758_U.if_write & AESL_inst_myproject.layer3_out_758_U.if_full_n;
    assign fifo_intf_2111.fifo_rd_block = 0;
    assign fifo_intf_2111.fifo_wr_block = 0;
    assign fifo_intf_2111.finish = finish;
    csv_file_dump fifo_csv_dumper_2111;
    csv_file_dump cstatus_csv_dumper_2111;
    df_fifo_monitor fifo_monitor_2111;
    df_fifo_intf fifo_intf_2112(clock,reset);
    assign fifo_intf_2112.rd_en = AESL_inst_myproject.layer3_out_759_U.if_read & AESL_inst_myproject.layer3_out_759_U.if_empty_n;
    assign fifo_intf_2112.wr_en = AESL_inst_myproject.layer3_out_759_U.if_write & AESL_inst_myproject.layer3_out_759_U.if_full_n;
    assign fifo_intf_2112.fifo_rd_block = 0;
    assign fifo_intf_2112.fifo_wr_block = 0;
    assign fifo_intf_2112.finish = finish;
    csv_file_dump fifo_csv_dumper_2112;
    csv_file_dump cstatus_csv_dumper_2112;
    df_fifo_monitor fifo_monitor_2112;
    df_fifo_intf fifo_intf_2113(clock,reset);
    assign fifo_intf_2113.rd_en = AESL_inst_myproject.layer3_out_760_U.if_read & AESL_inst_myproject.layer3_out_760_U.if_empty_n;
    assign fifo_intf_2113.wr_en = AESL_inst_myproject.layer3_out_760_U.if_write & AESL_inst_myproject.layer3_out_760_U.if_full_n;
    assign fifo_intf_2113.fifo_rd_block = 0;
    assign fifo_intf_2113.fifo_wr_block = 0;
    assign fifo_intf_2113.finish = finish;
    csv_file_dump fifo_csv_dumper_2113;
    csv_file_dump cstatus_csv_dumper_2113;
    df_fifo_monitor fifo_monitor_2113;
    df_fifo_intf fifo_intf_2114(clock,reset);
    assign fifo_intf_2114.rd_en = AESL_inst_myproject.layer3_out_761_U.if_read & AESL_inst_myproject.layer3_out_761_U.if_empty_n;
    assign fifo_intf_2114.wr_en = AESL_inst_myproject.layer3_out_761_U.if_write & AESL_inst_myproject.layer3_out_761_U.if_full_n;
    assign fifo_intf_2114.fifo_rd_block = 0;
    assign fifo_intf_2114.fifo_wr_block = 0;
    assign fifo_intf_2114.finish = finish;
    csv_file_dump fifo_csv_dumper_2114;
    csv_file_dump cstatus_csv_dumper_2114;
    df_fifo_monitor fifo_monitor_2114;
    df_fifo_intf fifo_intf_2115(clock,reset);
    assign fifo_intf_2115.rd_en = AESL_inst_myproject.layer3_out_762_U.if_read & AESL_inst_myproject.layer3_out_762_U.if_empty_n;
    assign fifo_intf_2115.wr_en = AESL_inst_myproject.layer3_out_762_U.if_write & AESL_inst_myproject.layer3_out_762_U.if_full_n;
    assign fifo_intf_2115.fifo_rd_block = 0;
    assign fifo_intf_2115.fifo_wr_block = 0;
    assign fifo_intf_2115.finish = finish;
    csv_file_dump fifo_csv_dumper_2115;
    csv_file_dump cstatus_csv_dumper_2115;
    df_fifo_monitor fifo_monitor_2115;
    df_fifo_intf fifo_intf_2116(clock,reset);
    assign fifo_intf_2116.rd_en = AESL_inst_myproject.layer3_out_763_U.if_read & AESL_inst_myproject.layer3_out_763_U.if_empty_n;
    assign fifo_intf_2116.wr_en = AESL_inst_myproject.layer3_out_763_U.if_write & AESL_inst_myproject.layer3_out_763_U.if_full_n;
    assign fifo_intf_2116.fifo_rd_block = 0;
    assign fifo_intf_2116.fifo_wr_block = 0;
    assign fifo_intf_2116.finish = finish;
    csv_file_dump fifo_csv_dumper_2116;
    csv_file_dump cstatus_csv_dumper_2116;
    df_fifo_monitor fifo_monitor_2116;
    df_fifo_intf fifo_intf_2117(clock,reset);
    assign fifo_intf_2117.rd_en = AESL_inst_myproject.layer3_out_764_U.if_read & AESL_inst_myproject.layer3_out_764_U.if_empty_n;
    assign fifo_intf_2117.wr_en = AESL_inst_myproject.layer3_out_764_U.if_write & AESL_inst_myproject.layer3_out_764_U.if_full_n;
    assign fifo_intf_2117.fifo_rd_block = 0;
    assign fifo_intf_2117.fifo_wr_block = 0;
    assign fifo_intf_2117.finish = finish;
    csv_file_dump fifo_csv_dumper_2117;
    csv_file_dump cstatus_csv_dumper_2117;
    df_fifo_monitor fifo_monitor_2117;
    df_fifo_intf fifo_intf_2118(clock,reset);
    assign fifo_intf_2118.rd_en = AESL_inst_myproject.layer3_out_765_U.if_read & AESL_inst_myproject.layer3_out_765_U.if_empty_n;
    assign fifo_intf_2118.wr_en = AESL_inst_myproject.layer3_out_765_U.if_write & AESL_inst_myproject.layer3_out_765_U.if_full_n;
    assign fifo_intf_2118.fifo_rd_block = 0;
    assign fifo_intf_2118.fifo_wr_block = 0;
    assign fifo_intf_2118.finish = finish;
    csv_file_dump fifo_csv_dumper_2118;
    csv_file_dump cstatus_csv_dumper_2118;
    df_fifo_monitor fifo_monitor_2118;
    df_fifo_intf fifo_intf_2119(clock,reset);
    assign fifo_intf_2119.rd_en = AESL_inst_myproject.layer3_out_766_U.if_read & AESL_inst_myproject.layer3_out_766_U.if_empty_n;
    assign fifo_intf_2119.wr_en = AESL_inst_myproject.layer3_out_766_U.if_write & AESL_inst_myproject.layer3_out_766_U.if_full_n;
    assign fifo_intf_2119.fifo_rd_block = 0;
    assign fifo_intf_2119.fifo_wr_block = 0;
    assign fifo_intf_2119.finish = finish;
    csv_file_dump fifo_csv_dumper_2119;
    csv_file_dump cstatus_csv_dumper_2119;
    df_fifo_monitor fifo_monitor_2119;
    df_fifo_intf fifo_intf_2120(clock,reset);
    assign fifo_intf_2120.rd_en = AESL_inst_myproject.layer3_out_767_U.if_read & AESL_inst_myproject.layer3_out_767_U.if_empty_n;
    assign fifo_intf_2120.wr_en = AESL_inst_myproject.layer3_out_767_U.if_write & AESL_inst_myproject.layer3_out_767_U.if_full_n;
    assign fifo_intf_2120.fifo_rd_block = 0;
    assign fifo_intf_2120.fifo_wr_block = 0;
    assign fifo_intf_2120.finish = finish;
    csv_file_dump fifo_csv_dumper_2120;
    csv_file_dump cstatus_csv_dumper_2120;
    df_fifo_monitor fifo_monitor_2120;
    df_fifo_intf fifo_intf_2121(clock,reset);
    assign fifo_intf_2121.rd_en = AESL_inst_myproject.layer3_out_768_U.if_read & AESL_inst_myproject.layer3_out_768_U.if_empty_n;
    assign fifo_intf_2121.wr_en = AESL_inst_myproject.layer3_out_768_U.if_write & AESL_inst_myproject.layer3_out_768_U.if_full_n;
    assign fifo_intf_2121.fifo_rd_block = 0;
    assign fifo_intf_2121.fifo_wr_block = 0;
    assign fifo_intf_2121.finish = finish;
    csv_file_dump fifo_csv_dumper_2121;
    csv_file_dump cstatus_csv_dumper_2121;
    df_fifo_monitor fifo_monitor_2121;
    df_fifo_intf fifo_intf_2122(clock,reset);
    assign fifo_intf_2122.rd_en = AESL_inst_myproject.layer3_out_769_U.if_read & AESL_inst_myproject.layer3_out_769_U.if_empty_n;
    assign fifo_intf_2122.wr_en = AESL_inst_myproject.layer3_out_769_U.if_write & AESL_inst_myproject.layer3_out_769_U.if_full_n;
    assign fifo_intf_2122.fifo_rd_block = 0;
    assign fifo_intf_2122.fifo_wr_block = 0;
    assign fifo_intf_2122.finish = finish;
    csv_file_dump fifo_csv_dumper_2122;
    csv_file_dump cstatus_csv_dumper_2122;
    df_fifo_monitor fifo_monitor_2122;
    df_fifo_intf fifo_intf_2123(clock,reset);
    assign fifo_intf_2123.rd_en = AESL_inst_myproject.layer3_out_770_U.if_read & AESL_inst_myproject.layer3_out_770_U.if_empty_n;
    assign fifo_intf_2123.wr_en = AESL_inst_myproject.layer3_out_770_U.if_write & AESL_inst_myproject.layer3_out_770_U.if_full_n;
    assign fifo_intf_2123.fifo_rd_block = 0;
    assign fifo_intf_2123.fifo_wr_block = 0;
    assign fifo_intf_2123.finish = finish;
    csv_file_dump fifo_csv_dumper_2123;
    csv_file_dump cstatus_csv_dumper_2123;
    df_fifo_monitor fifo_monitor_2123;
    df_fifo_intf fifo_intf_2124(clock,reset);
    assign fifo_intf_2124.rd_en = AESL_inst_myproject.layer3_out_771_U.if_read & AESL_inst_myproject.layer3_out_771_U.if_empty_n;
    assign fifo_intf_2124.wr_en = AESL_inst_myproject.layer3_out_771_U.if_write & AESL_inst_myproject.layer3_out_771_U.if_full_n;
    assign fifo_intf_2124.fifo_rd_block = 0;
    assign fifo_intf_2124.fifo_wr_block = 0;
    assign fifo_intf_2124.finish = finish;
    csv_file_dump fifo_csv_dumper_2124;
    csv_file_dump cstatus_csv_dumper_2124;
    df_fifo_monitor fifo_monitor_2124;
    df_fifo_intf fifo_intf_2125(clock,reset);
    assign fifo_intf_2125.rd_en = AESL_inst_myproject.layer3_out_772_U.if_read & AESL_inst_myproject.layer3_out_772_U.if_empty_n;
    assign fifo_intf_2125.wr_en = AESL_inst_myproject.layer3_out_772_U.if_write & AESL_inst_myproject.layer3_out_772_U.if_full_n;
    assign fifo_intf_2125.fifo_rd_block = 0;
    assign fifo_intf_2125.fifo_wr_block = 0;
    assign fifo_intf_2125.finish = finish;
    csv_file_dump fifo_csv_dumper_2125;
    csv_file_dump cstatus_csv_dumper_2125;
    df_fifo_monitor fifo_monitor_2125;
    df_fifo_intf fifo_intf_2126(clock,reset);
    assign fifo_intf_2126.rd_en = AESL_inst_myproject.layer3_out_773_U.if_read & AESL_inst_myproject.layer3_out_773_U.if_empty_n;
    assign fifo_intf_2126.wr_en = AESL_inst_myproject.layer3_out_773_U.if_write & AESL_inst_myproject.layer3_out_773_U.if_full_n;
    assign fifo_intf_2126.fifo_rd_block = 0;
    assign fifo_intf_2126.fifo_wr_block = 0;
    assign fifo_intf_2126.finish = finish;
    csv_file_dump fifo_csv_dumper_2126;
    csv_file_dump cstatus_csv_dumper_2126;
    df_fifo_monitor fifo_monitor_2126;
    df_fifo_intf fifo_intf_2127(clock,reset);
    assign fifo_intf_2127.rd_en = AESL_inst_myproject.layer3_out_774_U.if_read & AESL_inst_myproject.layer3_out_774_U.if_empty_n;
    assign fifo_intf_2127.wr_en = AESL_inst_myproject.layer3_out_774_U.if_write & AESL_inst_myproject.layer3_out_774_U.if_full_n;
    assign fifo_intf_2127.fifo_rd_block = 0;
    assign fifo_intf_2127.fifo_wr_block = 0;
    assign fifo_intf_2127.finish = finish;
    csv_file_dump fifo_csv_dumper_2127;
    csv_file_dump cstatus_csv_dumper_2127;
    df_fifo_monitor fifo_monitor_2127;
    df_fifo_intf fifo_intf_2128(clock,reset);
    assign fifo_intf_2128.rd_en = AESL_inst_myproject.layer3_out_775_U.if_read & AESL_inst_myproject.layer3_out_775_U.if_empty_n;
    assign fifo_intf_2128.wr_en = AESL_inst_myproject.layer3_out_775_U.if_write & AESL_inst_myproject.layer3_out_775_U.if_full_n;
    assign fifo_intf_2128.fifo_rd_block = 0;
    assign fifo_intf_2128.fifo_wr_block = 0;
    assign fifo_intf_2128.finish = finish;
    csv_file_dump fifo_csv_dumper_2128;
    csv_file_dump cstatus_csv_dumper_2128;
    df_fifo_monitor fifo_monitor_2128;
    df_fifo_intf fifo_intf_2129(clock,reset);
    assign fifo_intf_2129.rd_en = AESL_inst_myproject.layer3_out_776_U.if_read & AESL_inst_myproject.layer3_out_776_U.if_empty_n;
    assign fifo_intf_2129.wr_en = AESL_inst_myproject.layer3_out_776_U.if_write & AESL_inst_myproject.layer3_out_776_U.if_full_n;
    assign fifo_intf_2129.fifo_rd_block = 0;
    assign fifo_intf_2129.fifo_wr_block = 0;
    assign fifo_intf_2129.finish = finish;
    csv_file_dump fifo_csv_dumper_2129;
    csv_file_dump cstatus_csv_dumper_2129;
    df_fifo_monitor fifo_monitor_2129;
    df_fifo_intf fifo_intf_2130(clock,reset);
    assign fifo_intf_2130.rd_en = AESL_inst_myproject.layer3_out_777_U.if_read & AESL_inst_myproject.layer3_out_777_U.if_empty_n;
    assign fifo_intf_2130.wr_en = AESL_inst_myproject.layer3_out_777_U.if_write & AESL_inst_myproject.layer3_out_777_U.if_full_n;
    assign fifo_intf_2130.fifo_rd_block = 0;
    assign fifo_intf_2130.fifo_wr_block = 0;
    assign fifo_intf_2130.finish = finish;
    csv_file_dump fifo_csv_dumper_2130;
    csv_file_dump cstatus_csv_dumper_2130;
    df_fifo_monitor fifo_monitor_2130;
    df_fifo_intf fifo_intf_2131(clock,reset);
    assign fifo_intf_2131.rd_en = AESL_inst_myproject.layer3_out_778_U.if_read & AESL_inst_myproject.layer3_out_778_U.if_empty_n;
    assign fifo_intf_2131.wr_en = AESL_inst_myproject.layer3_out_778_U.if_write & AESL_inst_myproject.layer3_out_778_U.if_full_n;
    assign fifo_intf_2131.fifo_rd_block = 0;
    assign fifo_intf_2131.fifo_wr_block = 0;
    assign fifo_intf_2131.finish = finish;
    csv_file_dump fifo_csv_dumper_2131;
    csv_file_dump cstatus_csv_dumper_2131;
    df_fifo_monitor fifo_monitor_2131;
    df_fifo_intf fifo_intf_2132(clock,reset);
    assign fifo_intf_2132.rd_en = AESL_inst_myproject.layer3_out_779_U.if_read & AESL_inst_myproject.layer3_out_779_U.if_empty_n;
    assign fifo_intf_2132.wr_en = AESL_inst_myproject.layer3_out_779_U.if_write & AESL_inst_myproject.layer3_out_779_U.if_full_n;
    assign fifo_intf_2132.fifo_rd_block = 0;
    assign fifo_intf_2132.fifo_wr_block = 0;
    assign fifo_intf_2132.finish = finish;
    csv_file_dump fifo_csv_dumper_2132;
    csv_file_dump cstatus_csv_dumper_2132;
    df_fifo_monitor fifo_monitor_2132;
    df_fifo_intf fifo_intf_2133(clock,reset);
    assign fifo_intf_2133.rd_en = AESL_inst_myproject.layer3_out_780_U.if_read & AESL_inst_myproject.layer3_out_780_U.if_empty_n;
    assign fifo_intf_2133.wr_en = AESL_inst_myproject.layer3_out_780_U.if_write & AESL_inst_myproject.layer3_out_780_U.if_full_n;
    assign fifo_intf_2133.fifo_rd_block = 0;
    assign fifo_intf_2133.fifo_wr_block = 0;
    assign fifo_intf_2133.finish = finish;
    csv_file_dump fifo_csv_dumper_2133;
    csv_file_dump cstatus_csv_dumper_2133;
    df_fifo_monitor fifo_monitor_2133;
    df_fifo_intf fifo_intf_2134(clock,reset);
    assign fifo_intf_2134.rd_en = AESL_inst_myproject.layer3_out_781_U.if_read & AESL_inst_myproject.layer3_out_781_U.if_empty_n;
    assign fifo_intf_2134.wr_en = AESL_inst_myproject.layer3_out_781_U.if_write & AESL_inst_myproject.layer3_out_781_U.if_full_n;
    assign fifo_intf_2134.fifo_rd_block = 0;
    assign fifo_intf_2134.fifo_wr_block = 0;
    assign fifo_intf_2134.finish = finish;
    csv_file_dump fifo_csv_dumper_2134;
    csv_file_dump cstatus_csv_dumper_2134;
    df_fifo_monitor fifo_monitor_2134;
    df_fifo_intf fifo_intf_2135(clock,reset);
    assign fifo_intf_2135.rd_en = AESL_inst_myproject.layer3_out_782_U.if_read & AESL_inst_myproject.layer3_out_782_U.if_empty_n;
    assign fifo_intf_2135.wr_en = AESL_inst_myproject.layer3_out_782_U.if_write & AESL_inst_myproject.layer3_out_782_U.if_full_n;
    assign fifo_intf_2135.fifo_rd_block = 0;
    assign fifo_intf_2135.fifo_wr_block = 0;
    assign fifo_intf_2135.finish = finish;
    csv_file_dump fifo_csv_dumper_2135;
    csv_file_dump cstatus_csv_dumper_2135;
    df_fifo_monitor fifo_monitor_2135;
    df_fifo_intf fifo_intf_2136(clock,reset);
    assign fifo_intf_2136.rd_en = AESL_inst_myproject.layer3_out_783_U.if_read & AESL_inst_myproject.layer3_out_783_U.if_empty_n;
    assign fifo_intf_2136.wr_en = AESL_inst_myproject.layer3_out_783_U.if_write & AESL_inst_myproject.layer3_out_783_U.if_full_n;
    assign fifo_intf_2136.fifo_rd_block = 0;
    assign fifo_intf_2136.fifo_wr_block = 0;
    assign fifo_intf_2136.finish = finish;
    csv_file_dump fifo_csv_dumper_2136;
    csv_file_dump cstatus_csv_dumper_2136;
    df_fifo_monitor fifo_monitor_2136;
    df_fifo_intf fifo_intf_2137(clock,reset);
    assign fifo_intf_2137.rd_en = AESL_inst_myproject.layer3_out_784_U.if_read & AESL_inst_myproject.layer3_out_784_U.if_empty_n;
    assign fifo_intf_2137.wr_en = AESL_inst_myproject.layer3_out_784_U.if_write & AESL_inst_myproject.layer3_out_784_U.if_full_n;
    assign fifo_intf_2137.fifo_rd_block = 0;
    assign fifo_intf_2137.fifo_wr_block = 0;
    assign fifo_intf_2137.finish = finish;
    csv_file_dump fifo_csv_dumper_2137;
    csv_file_dump cstatus_csv_dumper_2137;
    df_fifo_monitor fifo_monitor_2137;
    df_fifo_intf fifo_intf_2138(clock,reset);
    assign fifo_intf_2138.rd_en = AESL_inst_myproject.layer3_out_785_U.if_read & AESL_inst_myproject.layer3_out_785_U.if_empty_n;
    assign fifo_intf_2138.wr_en = AESL_inst_myproject.layer3_out_785_U.if_write & AESL_inst_myproject.layer3_out_785_U.if_full_n;
    assign fifo_intf_2138.fifo_rd_block = 0;
    assign fifo_intf_2138.fifo_wr_block = 0;
    assign fifo_intf_2138.finish = finish;
    csv_file_dump fifo_csv_dumper_2138;
    csv_file_dump cstatus_csv_dumper_2138;
    df_fifo_monitor fifo_monitor_2138;
    df_fifo_intf fifo_intf_2139(clock,reset);
    assign fifo_intf_2139.rd_en = AESL_inst_myproject.layer3_out_786_U.if_read & AESL_inst_myproject.layer3_out_786_U.if_empty_n;
    assign fifo_intf_2139.wr_en = AESL_inst_myproject.layer3_out_786_U.if_write & AESL_inst_myproject.layer3_out_786_U.if_full_n;
    assign fifo_intf_2139.fifo_rd_block = 0;
    assign fifo_intf_2139.fifo_wr_block = 0;
    assign fifo_intf_2139.finish = finish;
    csv_file_dump fifo_csv_dumper_2139;
    csv_file_dump cstatus_csv_dumper_2139;
    df_fifo_monitor fifo_monitor_2139;
    df_fifo_intf fifo_intf_2140(clock,reset);
    assign fifo_intf_2140.rd_en = AESL_inst_myproject.layer3_out_787_U.if_read & AESL_inst_myproject.layer3_out_787_U.if_empty_n;
    assign fifo_intf_2140.wr_en = AESL_inst_myproject.layer3_out_787_U.if_write & AESL_inst_myproject.layer3_out_787_U.if_full_n;
    assign fifo_intf_2140.fifo_rd_block = 0;
    assign fifo_intf_2140.fifo_wr_block = 0;
    assign fifo_intf_2140.finish = finish;
    csv_file_dump fifo_csv_dumper_2140;
    csv_file_dump cstatus_csv_dumper_2140;
    df_fifo_monitor fifo_monitor_2140;
    df_fifo_intf fifo_intf_2141(clock,reset);
    assign fifo_intf_2141.rd_en = AESL_inst_myproject.layer3_out_788_U.if_read & AESL_inst_myproject.layer3_out_788_U.if_empty_n;
    assign fifo_intf_2141.wr_en = AESL_inst_myproject.layer3_out_788_U.if_write & AESL_inst_myproject.layer3_out_788_U.if_full_n;
    assign fifo_intf_2141.fifo_rd_block = 0;
    assign fifo_intf_2141.fifo_wr_block = 0;
    assign fifo_intf_2141.finish = finish;
    csv_file_dump fifo_csv_dumper_2141;
    csv_file_dump cstatus_csv_dumper_2141;
    df_fifo_monitor fifo_monitor_2141;
    df_fifo_intf fifo_intf_2142(clock,reset);
    assign fifo_intf_2142.rd_en = AESL_inst_myproject.layer3_out_789_U.if_read & AESL_inst_myproject.layer3_out_789_U.if_empty_n;
    assign fifo_intf_2142.wr_en = AESL_inst_myproject.layer3_out_789_U.if_write & AESL_inst_myproject.layer3_out_789_U.if_full_n;
    assign fifo_intf_2142.fifo_rd_block = 0;
    assign fifo_intf_2142.fifo_wr_block = 0;
    assign fifo_intf_2142.finish = finish;
    csv_file_dump fifo_csv_dumper_2142;
    csv_file_dump cstatus_csv_dumper_2142;
    df_fifo_monitor fifo_monitor_2142;
    df_fifo_intf fifo_intf_2143(clock,reset);
    assign fifo_intf_2143.rd_en = AESL_inst_myproject.layer3_out_790_U.if_read & AESL_inst_myproject.layer3_out_790_U.if_empty_n;
    assign fifo_intf_2143.wr_en = AESL_inst_myproject.layer3_out_790_U.if_write & AESL_inst_myproject.layer3_out_790_U.if_full_n;
    assign fifo_intf_2143.fifo_rd_block = 0;
    assign fifo_intf_2143.fifo_wr_block = 0;
    assign fifo_intf_2143.finish = finish;
    csv_file_dump fifo_csv_dumper_2143;
    csv_file_dump cstatus_csv_dumper_2143;
    df_fifo_monitor fifo_monitor_2143;
    df_fifo_intf fifo_intf_2144(clock,reset);
    assign fifo_intf_2144.rd_en = AESL_inst_myproject.layer3_out_791_U.if_read & AESL_inst_myproject.layer3_out_791_U.if_empty_n;
    assign fifo_intf_2144.wr_en = AESL_inst_myproject.layer3_out_791_U.if_write & AESL_inst_myproject.layer3_out_791_U.if_full_n;
    assign fifo_intf_2144.fifo_rd_block = 0;
    assign fifo_intf_2144.fifo_wr_block = 0;
    assign fifo_intf_2144.finish = finish;
    csv_file_dump fifo_csv_dumper_2144;
    csv_file_dump cstatus_csv_dumper_2144;
    df_fifo_monitor fifo_monitor_2144;
    df_fifo_intf fifo_intf_2145(clock,reset);
    assign fifo_intf_2145.rd_en = AESL_inst_myproject.layer3_out_792_U.if_read & AESL_inst_myproject.layer3_out_792_U.if_empty_n;
    assign fifo_intf_2145.wr_en = AESL_inst_myproject.layer3_out_792_U.if_write & AESL_inst_myproject.layer3_out_792_U.if_full_n;
    assign fifo_intf_2145.fifo_rd_block = 0;
    assign fifo_intf_2145.fifo_wr_block = 0;
    assign fifo_intf_2145.finish = finish;
    csv_file_dump fifo_csv_dumper_2145;
    csv_file_dump cstatus_csv_dumper_2145;
    df_fifo_monitor fifo_monitor_2145;
    df_fifo_intf fifo_intf_2146(clock,reset);
    assign fifo_intf_2146.rd_en = AESL_inst_myproject.layer3_out_793_U.if_read & AESL_inst_myproject.layer3_out_793_U.if_empty_n;
    assign fifo_intf_2146.wr_en = AESL_inst_myproject.layer3_out_793_U.if_write & AESL_inst_myproject.layer3_out_793_U.if_full_n;
    assign fifo_intf_2146.fifo_rd_block = 0;
    assign fifo_intf_2146.fifo_wr_block = 0;
    assign fifo_intf_2146.finish = finish;
    csv_file_dump fifo_csv_dumper_2146;
    csv_file_dump cstatus_csv_dumper_2146;
    df_fifo_monitor fifo_monitor_2146;
    df_fifo_intf fifo_intf_2147(clock,reset);
    assign fifo_intf_2147.rd_en = AESL_inst_myproject.layer3_out_794_U.if_read & AESL_inst_myproject.layer3_out_794_U.if_empty_n;
    assign fifo_intf_2147.wr_en = AESL_inst_myproject.layer3_out_794_U.if_write & AESL_inst_myproject.layer3_out_794_U.if_full_n;
    assign fifo_intf_2147.fifo_rd_block = 0;
    assign fifo_intf_2147.fifo_wr_block = 0;
    assign fifo_intf_2147.finish = finish;
    csv_file_dump fifo_csv_dumper_2147;
    csv_file_dump cstatus_csv_dumper_2147;
    df_fifo_monitor fifo_monitor_2147;
    df_fifo_intf fifo_intf_2148(clock,reset);
    assign fifo_intf_2148.rd_en = AESL_inst_myproject.layer3_out_795_U.if_read & AESL_inst_myproject.layer3_out_795_U.if_empty_n;
    assign fifo_intf_2148.wr_en = AESL_inst_myproject.layer3_out_795_U.if_write & AESL_inst_myproject.layer3_out_795_U.if_full_n;
    assign fifo_intf_2148.fifo_rd_block = 0;
    assign fifo_intf_2148.fifo_wr_block = 0;
    assign fifo_intf_2148.finish = finish;
    csv_file_dump fifo_csv_dumper_2148;
    csv_file_dump cstatus_csv_dumper_2148;
    df_fifo_monitor fifo_monitor_2148;
    df_fifo_intf fifo_intf_2149(clock,reset);
    assign fifo_intf_2149.rd_en = AESL_inst_myproject.layer3_out_796_U.if_read & AESL_inst_myproject.layer3_out_796_U.if_empty_n;
    assign fifo_intf_2149.wr_en = AESL_inst_myproject.layer3_out_796_U.if_write & AESL_inst_myproject.layer3_out_796_U.if_full_n;
    assign fifo_intf_2149.fifo_rd_block = 0;
    assign fifo_intf_2149.fifo_wr_block = 0;
    assign fifo_intf_2149.finish = finish;
    csv_file_dump fifo_csv_dumper_2149;
    csv_file_dump cstatus_csv_dumper_2149;
    df_fifo_monitor fifo_monitor_2149;
    df_fifo_intf fifo_intf_2150(clock,reset);
    assign fifo_intf_2150.rd_en = AESL_inst_myproject.layer3_out_797_U.if_read & AESL_inst_myproject.layer3_out_797_U.if_empty_n;
    assign fifo_intf_2150.wr_en = AESL_inst_myproject.layer3_out_797_U.if_write & AESL_inst_myproject.layer3_out_797_U.if_full_n;
    assign fifo_intf_2150.fifo_rd_block = 0;
    assign fifo_intf_2150.fifo_wr_block = 0;
    assign fifo_intf_2150.finish = finish;
    csv_file_dump fifo_csv_dumper_2150;
    csv_file_dump cstatus_csv_dumper_2150;
    df_fifo_monitor fifo_monitor_2150;
    df_fifo_intf fifo_intf_2151(clock,reset);
    assign fifo_intf_2151.rd_en = AESL_inst_myproject.layer3_out_798_U.if_read & AESL_inst_myproject.layer3_out_798_U.if_empty_n;
    assign fifo_intf_2151.wr_en = AESL_inst_myproject.layer3_out_798_U.if_write & AESL_inst_myproject.layer3_out_798_U.if_full_n;
    assign fifo_intf_2151.fifo_rd_block = 0;
    assign fifo_intf_2151.fifo_wr_block = 0;
    assign fifo_intf_2151.finish = finish;
    csv_file_dump fifo_csv_dumper_2151;
    csv_file_dump cstatus_csv_dumper_2151;
    df_fifo_monitor fifo_monitor_2151;
    df_fifo_intf fifo_intf_2152(clock,reset);
    assign fifo_intf_2152.rd_en = AESL_inst_myproject.layer3_out_799_U.if_read & AESL_inst_myproject.layer3_out_799_U.if_empty_n;
    assign fifo_intf_2152.wr_en = AESL_inst_myproject.layer3_out_799_U.if_write & AESL_inst_myproject.layer3_out_799_U.if_full_n;
    assign fifo_intf_2152.fifo_rd_block = 0;
    assign fifo_intf_2152.fifo_wr_block = 0;
    assign fifo_intf_2152.finish = finish;
    csv_file_dump fifo_csv_dumper_2152;
    csv_file_dump cstatus_csv_dumper_2152;
    df_fifo_monitor fifo_monitor_2152;
    df_fifo_intf fifo_intf_2153(clock,reset);
    assign fifo_intf_2153.rd_en = AESL_inst_myproject.layer3_out_800_U.if_read & AESL_inst_myproject.layer3_out_800_U.if_empty_n;
    assign fifo_intf_2153.wr_en = AESL_inst_myproject.layer3_out_800_U.if_write & AESL_inst_myproject.layer3_out_800_U.if_full_n;
    assign fifo_intf_2153.fifo_rd_block = 0;
    assign fifo_intf_2153.fifo_wr_block = 0;
    assign fifo_intf_2153.finish = finish;
    csv_file_dump fifo_csv_dumper_2153;
    csv_file_dump cstatus_csv_dumper_2153;
    df_fifo_monitor fifo_monitor_2153;
    df_fifo_intf fifo_intf_2154(clock,reset);
    assign fifo_intf_2154.rd_en = AESL_inst_myproject.layer3_out_801_U.if_read & AESL_inst_myproject.layer3_out_801_U.if_empty_n;
    assign fifo_intf_2154.wr_en = AESL_inst_myproject.layer3_out_801_U.if_write & AESL_inst_myproject.layer3_out_801_U.if_full_n;
    assign fifo_intf_2154.fifo_rd_block = 0;
    assign fifo_intf_2154.fifo_wr_block = 0;
    assign fifo_intf_2154.finish = finish;
    csv_file_dump fifo_csv_dumper_2154;
    csv_file_dump cstatus_csv_dumper_2154;
    df_fifo_monitor fifo_monitor_2154;
    df_fifo_intf fifo_intf_2155(clock,reset);
    assign fifo_intf_2155.rd_en = AESL_inst_myproject.layer3_out_802_U.if_read & AESL_inst_myproject.layer3_out_802_U.if_empty_n;
    assign fifo_intf_2155.wr_en = AESL_inst_myproject.layer3_out_802_U.if_write & AESL_inst_myproject.layer3_out_802_U.if_full_n;
    assign fifo_intf_2155.fifo_rd_block = 0;
    assign fifo_intf_2155.fifo_wr_block = 0;
    assign fifo_intf_2155.finish = finish;
    csv_file_dump fifo_csv_dumper_2155;
    csv_file_dump cstatus_csv_dumper_2155;
    df_fifo_monitor fifo_monitor_2155;
    df_fifo_intf fifo_intf_2156(clock,reset);
    assign fifo_intf_2156.rd_en = AESL_inst_myproject.layer3_out_803_U.if_read & AESL_inst_myproject.layer3_out_803_U.if_empty_n;
    assign fifo_intf_2156.wr_en = AESL_inst_myproject.layer3_out_803_U.if_write & AESL_inst_myproject.layer3_out_803_U.if_full_n;
    assign fifo_intf_2156.fifo_rd_block = 0;
    assign fifo_intf_2156.fifo_wr_block = 0;
    assign fifo_intf_2156.finish = finish;
    csv_file_dump fifo_csv_dumper_2156;
    csv_file_dump cstatus_csv_dumper_2156;
    df_fifo_monitor fifo_monitor_2156;
    df_fifo_intf fifo_intf_2157(clock,reset);
    assign fifo_intf_2157.rd_en = AESL_inst_myproject.layer3_out_804_U.if_read & AESL_inst_myproject.layer3_out_804_U.if_empty_n;
    assign fifo_intf_2157.wr_en = AESL_inst_myproject.layer3_out_804_U.if_write & AESL_inst_myproject.layer3_out_804_U.if_full_n;
    assign fifo_intf_2157.fifo_rd_block = 0;
    assign fifo_intf_2157.fifo_wr_block = 0;
    assign fifo_intf_2157.finish = finish;
    csv_file_dump fifo_csv_dumper_2157;
    csv_file_dump cstatus_csv_dumper_2157;
    df_fifo_monitor fifo_monitor_2157;
    df_fifo_intf fifo_intf_2158(clock,reset);
    assign fifo_intf_2158.rd_en = AESL_inst_myproject.layer3_out_805_U.if_read & AESL_inst_myproject.layer3_out_805_U.if_empty_n;
    assign fifo_intf_2158.wr_en = AESL_inst_myproject.layer3_out_805_U.if_write & AESL_inst_myproject.layer3_out_805_U.if_full_n;
    assign fifo_intf_2158.fifo_rd_block = 0;
    assign fifo_intf_2158.fifo_wr_block = 0;
    assign fifo_intf_2158.finish = finish;
    csv_file_dump fifo_csv_dumper_2158;
    csv_file_dump cstatus_csv_dumper_2158;
    df_fifo_monitor fifo_monitor_2158;
    df_fifo_intf fifo_intf_2159(clock,reset);
    assign fifo_intf_2159.rd_en = AESL_inst_myproject.layer3_out_806_U.if_read & AESL_inst_myproject.layer3_out_806_U.if_empty_n;
    assign fifo_intf_2159.wr_en = AESL_inst_myproject.layer3_out_806_U.if_write & AESL_inst_myproject.layer3_out_806_U.if_full_n;
    assign fifo_intf_2159.fifo_rd_block = 0;
    assign fifo_intf_2159.fifo_wr_block = 0;
    assign fifo_intf_2159.finish = finish;
    csv_file_dump fifo_csv_dumper_2159;
    csv_file_dump cstatus_csv_dumper_2159;
    df_fifo_monitor fifo_monitor_2159;
    df_fifo_intf fifo_intf_2160(clock,reset);
    assign fifo_intf_2160.rd_en = AESL_inst_myproject.layer3_out_807_U.if_read & AESL_inst_myproject.layer3_out_807_U.if_empty_n;
    assign fifo_intf_2160.wr_en = AESL_inst_myproject.layer3_out_807_U.if_write & AESL_inst_myproject.layer3_out_807_U.if_full_n;
    assign fifo_intf_2160.fifo_rd_block = 0;
    assign fifo_intf_2160.fifo_wr_block = 0;
    assign fifo_intf_2160.finish = finish;
    csv_file_dump fifo_csv_dumper_2160;
    csv_file_dump cstatus_csv_dumper_2160;
    df_fifo_monitor fifo_monitor_2160;
    df_fifo_intf fifo_intf_2161(clock,reset);
    assign fifo_intf_2161.rd_en = AESL_inst_myproject.layer3_out_808_U.if_read & AESL_inst_myproject.layer3_out_808_U.if_empty_n;
    assign fifo_intf_2161.wr_en = AESL_inst_myproject.layer3_out_808_U.if_write & AESL_inst_myproject.layer3_out_808_U.if_full_n;
    assign fifo_intf_2161.fifo_rd_block = 0;
    assign fifo_intf_2161.fifo_wr_block = 0;
    assign fifo_intf_2161.finish = finish;
    csv_file_dump fifo_csv_dumper_2161;
    csv_file_dump cstatus_csv_dumper_2161;
    df_fifo_monitor fifo_monitor_2161;
    df_fifo_intf fifo_intf_2162(clock,reset);
    assign fifo_intf_2162.rd_en = AESL_inst_myproject.layer3_out_809_U.if_read & AESL_inst_myproject.layer3_out_809_U.if_empty_n;
    assign fifo_intf_2162.wr_en = AESL_inst_myproject.layer3_out_809_U.if_write & AESL_inst_myproject.layer3_out_809_U.if_full_n;
    assign fifo_intf_2162.fifo_rd_block = 0;
    assign fifo_intf_2162.fifo_wr_block = 0;
    assign fifo_intf_2162.finish = finish;
    csv_file_dump fifo_csv_dumper_2162;
    csv_file_dump cstatus_csv_dumper_2162;
    df_fifo_monitor fifo_monitor_2162;
    df_fifo_intf fifo_intf_2163(clock,reset);
    assign fifo_intf_2163.rd_en = AESL_inst_myproject.layer3_out_810_U.if_read & AESL_inst_myproject.layer3_out_810_U.if_empty_n;
    assign fifo_intf_2163.wr_en = AESL_inst_myproject.layer3_out_810_U.if_write & AESL_inst_myproject.layer3_out_810_U.if_full_n;
    assign fifo_intf_2163.fifo_rd_block = 0;
    assign fifo_intf_2163.fifo_wr_block = 0;
    assign fifo_intf_2163.finish = finish;
    csv_file_dump fifo_csv_dumper_2163;
    csv_file_dump cstatus_csv_dumper_2163;
    df_fifo_monitor fifo_monitor_2163;
    df_fifo_intf fifo_intf_2164(clock,reset);
    assign fifo_intf_2164.rd_en = AESL_inst_myproject.layer3_out_811_U.if_read & AESL_inst_myproject.layer3_out_811_U.if_empty_n;
    assign fifo_intf_2164.wr_en = AESL_inst_myproject.layer3_out_811_U.if_write & AESL_inst_myproject.layer3_out_811_U.if_full_n;
    assign fifo_intf_2164.fifo_rd_block = 0;
    assign fifo_intf_2164.fifo_wr_block = 0;
    assign fifo_intf_2164.finish = finish;
    csv_file_dump fifo_csv_dumper_2164;
    csv_file_dump cstatus_csv_dumper_2164;
    df_fifo_monitor fifo_monitor_2164;
    df_fifo_intf fifo_intf_2165(clock,reset);
    assign fifo_intf_2165.rd_en = AESL_inst_myproject.layer3_out_812_U.if_read & AESL_inst_myproject.layer3_out_812_U.if_empty_n;
    assign fifo_intf_2165.wr_en = AESL_inst_myproject.layer3_out_812_U.if_write & AESL_inst_myproject.layer3_out_812_U.if_full_n;
    assign fifo_intf_2165.fifo_rd_block = 0;
    assign fifo_intf_2165.fifo_wr_block = 0;
    assign fifo_intf_2165.finish = finish;
    csv_file_dump fifo_csv_dumper_2165;
    csv_file_dump cstatus_csv_dumper_2165;
    df_fifo_monitor fifo_monitor_2165;
    df_fifo_intf fifo_intf_2166(clock,reset);
    assign fifo_intf_2166.rd_en = AESL_inst_myproject.layer3_out_813_U.if_read & AESL_inst_myproject.layer3_out_813_U.if_empty_n;
    assign fifo_intf_2166.wr_en = AESL_inst_myproject.layer3_out_813_U.if_write & AESL_inst_myproject.layer3_out_813_U.if_full_n;
    assign fifo_intf_2166.fifo_rd_block = 0;
    assign fifo_intf_2166.fifo_wr_block = 0;
    assign fifo_intf_2166.finish = finish;
    csv_file_dump fifo_csv_dumper_2166;
    csv_file_dump cstatus_csv_dumper_2166;
    df_fifo_monitor fifo_monitor_2166;
    df_fifo_intf fifo_intf_2167(clock,reset);
    assign fifo_intf_2167.rd_en = AESL_inst_myproject.layer3_out_814_U.if_read & AESL_inst_myproject.layer3_out_814_U.if_empty_n;
    assign fifo_intf_2167.wr_en = AESL_inst_myproject.layer3_out_814_U.if_write & AESL_inst_myproject.layer3_out_814_U.if_full_n;
    assign fifo_intf_2167.fifo_rd_block = 0;
    assign fifo_intf_2167.fifo_wr_block = 0;
    assign fifo_intf_2167.finish = finish;
    csv_file_dump fifo_csv_dumper_2167;
    csv_file_dump cstatus_csv_dumper_2167;
    df_fifo_monitor fifo_monitor_2167;
    df_fifo_intf fifo_intf_2168(clock,reset);
    assign fifo_intf_2168.rd_en = AESL_inst_myproject.layer3_out_815_U.if_read & AESL_inst_myproject.layer3_out_815_U.if_empty_n;
    assign fifo_intf_2168.wr_en = AESL_inst_myproject.layer3_out_815_U.if_write & AESL_inst_myproject.layer3_out_815_U.if_full_n;
    assign fifo_intf_2168.fifo_rd_block = 0;
    assign fifo_intf_2168.fifo_wr_block = 0;
    assign fifo_intf_2168.finish = finish;
    csv_file_dump fifo_csv_dumper_2168;
    csv_file_dump cstatus_csv_dumper_2168;
    df_fifo_monitor fifo_monitor_2168;
    df_fifo_intf fifo_intf_2169(clock,reset);
    assign fifo_intf_2169.rd_en = AESL_inst_myproject.layer3_out_816_U.if_read & AESL_inst_myproject.layer3_out_816_U.if_empty_n;
    assign fifo_intf_2169.wr_en = AESL_inst_myproject.layer3_out_816_U.if_write & AESL_inst_myproject.layer3_out_816_U.if_full_n;
    assign fifo_intf_2169.fifo_rd_block = 0;
    assign fifo_intf_2169.fifo_wr_block = 0;
    assign fifo_intf_2169.finish = finish;
    csv_file_dump fifo_csv_dumper_2169;
    csv_file_dump cstatus_csv_dumper_2169;
    df_fifo_monitor fifo_monitor_2169;
    df_fifo_intf fifo_intf_2170(clock,reset);
    assign fifo_intf_2170.rd_en = AESL_inst_myproject.layer3_out_817_U.if_read & AESL_inst_myproject.layer3_out_817_U.if_empty_n;
    assign fifo_intf_2170.wr_en = AESL_inst_myproject.layer3_out_817_U.if_write & AESL_inst_myproject.layer3_out_817_U.if_full_n;
    assign fifo_intf_2170.fifo_rd_block = 0;
    assign fifo_intf_2170.fifo_wr_block = 0;
    assign fifo_intf_2170.finish = finish;
    csv_file_dump fifo_csv_dumper_2170;
    csv_file_dump cstatus_csv_dumper_2170;
    df_fifo_monitor fifo_monitor_2170;
    df_fifo_intf fifo_intf_2171(clock,reset);
    assign fifo_intf_2171.rd_en = AESL_inst_myproject.layer3_out_818_U.if_read & AESL_inst_myproject.layer3_out_818_U.if_empty_n;
    assign fifo_intf_2171.wr_en = AESL_inst_myproject.layer3_out_818_U.if_write & AESL_inst_myproject.layer3_out_818_U.if_full_n;
    assign fifo_intf_2171.fifo_rd_block = 0;
    assign fifo_intf_2171.fifo_wr_block = 0;
    assign fifo_intf_2171.finish = finish;
    csv_file_dump fifo_csv_dumper_2171;
    csv_file_dump cstatus_csv_dumper_2171;
    df_fifo_monitor fifo_monitor_2171;
    df_fifo_intf fifo_intf_2172(clock,reset);
    assign fifo_intf_2172.rd_en = AESL_inst_myproject.layer3_out_819_U.if_read & AESL_inst_myproject.layer3_out_819_U.if_empty_n;
    assign fifo_intf_2172.wr_en = AESL_inst_myproject.layer3_out_819_U.if_write & AESL_inst_myproject.layer3_out_819_U.if_full_n;
    assign fifo_intf_2172.fifo_rd_block = 0;
    assign fifo_intf_2172.fifo_wr_block = 0;
    assign fifo_intf_2172.finish = finish;
    csv_file_dump fifo_csv_dumper_2172;
    csv_file_dump cstatus_csv_dumper_2172;
    df_fifo_monitor fifo_monitor_2172;
    df_fifo_intf fifo_intf_2173(clock,reset);
    assign fifo_intf_2173.rd_en = AESL_inst_myproject.layer3_out_820_U.if_read & AESL_inst_myproject.layer3_out_820_U.if_empty_n;
    assign fifo_intf_2173.wr_en = AESL_inst_myproject.layer3_out_820_U.if_write & AESL_inst_myproject.layer3_out_820_U.if_full_n;
    assign fifo_intf_2173.fifo_rd_block = 0;
    assign fifo_intf_2173.fifo_wr_block = 0;
    assign fifo_intf_2173.finish = finish;
    csv_file_dump fifo_csv_dumper_2173;
    csv_file_dump cstatus_csv_dumper_2173;
    df_fifo_monitor fifo_monitor_2173;
    df_fifo_intf fifo_intf_2174(clock,reset);
    assign fifo_intf_2174.rd_en = AESL_inst_myproject.layer3_out_821_U.if_read & AESL_inst_myproject.layer3_out_821_U.if_empty_n;
    assign fifo_intf_2174.wr_en = AESL_inst_myproject.layer3_out_821_U.if_write & AESL_inst_myproject.layer3_out_821_U.if_full_n;
    assign fifo_intf_2174.fifo_rd_block = 0;
    assign fifo_intf_2174.fifo_wr_block = 0;
    assign fifo_intf_2174.finish = finish;
    csv_file_dump fifo_csv_dumper_2174;
    csv_file_dump cstatus_csv_dumper_2174;
    df_fifo_monitor fifo_monitor_2174;
    df_fifo_intf fifo_intf_2175(clock,reset);
    assign fifo_intf_2175.rd_en = AESL_inst_myproject.layer3_out_822_U.if_read & AESL_inst_myproject.layer3_out_822_U.if_empty_n;
    assign fifo_intf_2175.wr_en = AESL_inst_myproject.layer3_out_822_U.if_write & AESL_inst_myproject.layer3_out_822_U.if_full_n;
    assign fifo_intf_2175.fifo_rd_block = 0;
    assign fifo_intf_2175.fifo_wr_block = 0;
    assign fifo_intf_2175.finish = finish;
    csv_file_dump fifo_csv_dumper_2175;
    csv_file_dump cstatus_csv_dumper_2175;
    df_fifo_monitor fifo_monitor_2175;
    df_fifo_intf fifo_intf_2176(clock,reset);
    assign fifo_intf_2176.rd_en = AESL_inst_myproject.layer3_out_823_U.if_read & AESL_inst_myproject.layer3_out_823_U.if_empty_n;
    assign fifo_intf_2176.wr_en = AESL_inst_myproject.layer3_out_823_U.if_write & AESL_inst_myproject.layer3_out_823_U.if_full_n;
    assign fifo_intf_2176.fifo_rd_block = 0;
    assign fifo_intf_2176.fifo_wr_block = 0;
    assign fifo_intf_2176.finish = finish;
    csv_file_dump fifo_csv_dumper_2176;
    csv_file_dump cstatus_csv_dumper_2176;
    df_fifo_monitor fifo_monitor_2176;
    df_fifo_intf fifo_intf_2177(clock,reset);
    assign fifo_intf_2177.rd_en = AESL_inst_myproject.layer3_out_824_U.if_read & AESL_inst_myproject.layer3_out_824_U.if_empty_n;
    assign fifo_intf_2177.wr_en = AESL_inst_myproject.layer3_out_824_U.if_write & AESL_inst_myproject.layer3_out_824_U.if_full_n;
    assign fifo_intf_2177.fifo_rd_block = 0;
    assign fifo_intf_2177.fifo_wr_block = 0;
    assign fifo_intf_2177.finish = finish;
    csv_file_dump fifo_csv_dumper_2177;
    csv_file_dump cstatus_csv_dumper_2177;
    df_fifo_monitor fifo_monitor_2177;
    df_fifo_intf fifo_intf_2178(clock,reset);
    assign fifo_intf_2178.rd_en = AESL_inst_myproject.layer3_out_825_U.if_read & AESL_inst_myproject.layer3_out_825_U.if_empty_n;
    assign fifo_intf_2178.wr_en = AESL_inst_myproject.layer3_out_825_U.if_write & AESL_inst_myproject.layer3_out_825_U.if_full_n;
    assign fifo_intf_2178.fifo_rd_block = 0;
    assign fifo_intf_2178.fifo_wr_block = 0;
    assign fifo_intf_2178.finish = finish;
    csv_file_dump fifo_csv_dumper_2178;
    csv_file_dump cstatus_csv_dumper_2178;
    df_fifo_monitor fifo_monitor_2178;
    df_fifo_intf fifo_intf_2179(clock,reset);
    assign fifo_intf_2179.rd_en = AESL_inst_myproject.layer3_out_826_U.if_read & AESL_inst_myproject.layer3_out_826_U.if_empty_n;
    assign fifo_intf_2179.wr_en = AESL_inst_myproject.layer3_out_826_U.if_write & AESL_inst_myproject.layer3_out_826_U.if_full_n;
    assign fifo_intf_2179.fifo_rd_block = 0;
    assign fifo_intf_2179.fifo_wr_block = 0;
    assign fifo_intf_2179.finish = finish;
    csv_file_dump fifo_csv_dumper_2179;
    csv_file_dump cstatus_csv_dumper_2179;
    df_fifo_monitor fifo_monitor_2179;
    df_fifo_intf fifo_intf_2180(clock,reset);
    assign fifo_intf_2180.rd_en = AESL_inst_myproject.layer3_out_827_U.if_read & AESL_inst_myproject.layer3_out_827_U.if_empty_n;
    assign fifo_intf_2180.wr_en = AESL_inst_myproject.layer3_out_827_U.if_write & AESL_inst_myproject.layer3_out_827_U.if_full_n;
    assign fifo_intf_2180.fifo_rd_block = 0;
    assign fifo_intf_2180.fifo_wr_block = 0;
    assign fifo_intf_2180.finish = finish;
    csv_file_dump fifo_csv_dumper_2180;
    csv_file_dump cstatus_csv_dumper_2180;
    df_fifo_monitor fifo_monitor_2180;
    df_fifo_intf fifo_intf_2181(clock,reset);
    assign fifo_intf_2181.rd_en = AESL_inst_myproject.layer3_out_828_U.if_read & AESL_inst_myproject.layer3_out_828_U.if_empty_n;
    assign fifo_intf_2181.wr_en = AESL_inst_myproject.layer3_out_828_U.if_write & AESL_inst_myproject.layer3_out_828_U.if_full_n;
    assign fifo_intf_2181.fifo_rd_block = 0;
    assign fifo_intf_2181.fifo_wr_block = 0;
    assign fifo_intf_2181.finish = finish;
    csv_file_dump fifo_csv_dumper_2181;
    csv_file_dump cstatus_csv_dumper_2181;
    df_fifo_monitor fifo_monitor_2181;
    df_fifo_intf fifo_intf_2182(clock,reset);
    assign fifo_intf_2182.rd_en = AESL_inst_myproject.layer3_out_829_U.if_read & AESL_inst_myproject.layer3_out_829_U.if_empty_n;
    assign fifo_intf_2182.wr_en = AESL_inst_myproject.layer3_out_829_U.if_write & AESL_inst_myproject.layer3_out_829_U.if_full_n;
    assign fifo_intf_2182.fifo_rd_block = 0;
    assign fifo_intf_2182.fifo_wr_block = 0;
    assign fifo_intf_2182.finish = finish;
    csv_file_dump fifo_csv_dumper_2182;
    csv_file_dump cstatus_csv_dumper_2182;
    df_fifo_monitor fifo_monitor_2182;
    df_fifo_intf fifo_intf_2183(clock,reset);
    assign fifo_intf_2183.rd_en = AESL_inst_myproject.layer3_out_830_U.if_read & AESL_inst_myproject.layer3_out_830_U.if_empty_n;
    assign fifo_intf_2183.wr_en = AESL_inst_myproject.layer3_out_830_U.if_write & AESL_inst_myproject.layer3_out_830_U.if_full_n;
    assign fifo_intf_2183.fifo_rd_block = 0;
    assign fifo_intf_2183.fifo_wr_block = 0;
    assign fifo_intf_2183.finish = finish;
    csv_file_dump fifo_csv_dumper_2183;
    csv_file_dump cstatus_csv_dumper_2183;
    df_fifo_monitor fifo_monitor_2183;
    df_fifo_intf fifo_intf_2184(clock,reset);
    assign fifo_intf_2184.rd_en = AESL_inst_myproject.layer3_out_831_U.if_read & AESL_inst_myproject.layer3_out_831_U.if_empty_n;
    assign fifo_intf_2184.wr_en = AESL_inst_myproject.layer3_out_831_U.if_write & AESL_inst_myproject.layer3_out_831_U.if_full_n;
    assign fifo_intf_2184.fifo_rd_block = 0;
    assign fifo_intf_2184.fifo_wr_block = 0;
    assign fifo_intf_2184.finish = finish;
    csv_file_dump fifo_csv_dumper_2184;
    csv_file_dump cstatus_csv_dumper_2184;
    df_fifo_monitor fifo_monitor_2184;
    df_fifo_intf fifo_intf_2185(clock,reset);
    assign fifo_intf_2185.rd_en = AESL_inst_myproject.layer3_out_832_U.if_read & AESL_inst_myproject.layer3_out_832_U.if_empty_n;
    assign fifo_intf_2185.wr_en = AESL_inst_myproject.layer3_out_832_U.if_write & AESL_inst_myproject.layer3_out_832_U.if_full_n;
    assign fifo_intf_2185.fifo_rd_block = 0;
    assign fifo_intf_2185.fifo_wr_block = 0;
    assign fifo_intf_2185.finish = finish;
    csv_file_dump fifo_csv_dumper_2185;
    csv_file_dump cstatus_csv_dumper_2185;
    df_fifo_monitor fifo_monitor_2185;
    df_fifo_intf fifo_intf_2186(clock,reset);
    assign fifo_intf_2186.rd_en = AESL_inst_myproject.layer3_out_833_U.if_read & AESL_inst_myproject.layer3_out_833_U.if_empty_n;
    assign fifo_intf_2186.wr_en = AESL_inst_myproject.layer3_out_833_U.if_write & AESL_inst_myproject.layer3_out_833_U.if_full_n;
    assign fifo_intf_2186.fifo_rd_block = 0;
    assign fifo_intf_2186.fifo_wr_block = 0;
    assign fifo_intf_2186.finish = finish;
    csv_file_dump fifo_csv_dumper_2186;
    csv_file_dump cstatus_csv_dumper_2186;
    df_fifo_monitor fifo_monitor_2186;
    df_fifo_intf fifo_intf_2187(clock,reset);
    assign fifo_intf_2187.rd_en = AESL_inst_myproject.layer3_out_834_U.if_read & AESL_inst_myproject.layer3_out_834_U.if_empty_n;
    assign fifo_intf_2187.wr_en = AESL_inst_myproject.layer3_out_834_U.if_write & AESL_inst_myproject.layer3_out_834_U.if_full_n;
    assign fifo_intf_2187.fifo_rd_block = 0;
    assign fifo_intf_2187.fifo_wr_block = 0;
    assign fifo_intf_2187.finish = finish;
    csv_file_dump fifo_csv_dumper_2187;
    csv_file_dump cstatus_csv_dumper_2187;
    df_fifo_monitor fifo_monitor_2187;
    df_fifo_intf fifo_intf_2188(clock,reset);
    assign fifo_intf_2188.rd_en = AESL_inst_myproject.layer3_out_835_U.if_read & AESL_inst_myproject.layer3_out_835_U.if_empty_n;
    assign fifo_intf_2188.wr_en = AESL_inst_myproject.layer3_out_835_U.if_write & AESL_inst_myproject.layer3_out_835_U.if_full_n;
    assign fifo_intf_2188.fifo_rd_block = 0;
    assign fifo_intf_2188.fifo_wr_block = 0;
    assign fifo_intf_2188.finish = finish;
    csv_file_dump fifo_csv_dumper_2188;
    csv_file_dump cstatus_csv_dumper_2188;
    df_fifo_monitor fifo_monitor_2188;
    df_fifo_intf fifo_intf_2189(clock,reset);
    assign fifo_intf_2189.rd_en = AESL_inst_myproject.layer3_out_836_U.if_read & AESL_inst_myproject.layer3_out_836_U.if_empty_n;
    assign fifo_intf_2189.wr_en = AESL_inst_myproject.layer3_out_836_U.if_write & AESL_inst_myproject.layer3_out_836_U.if_full_n;
    assign fifo_intf_2189.fifo_rd_block = 0;
    assign fifo_intf_2189.fifo_wr_block = 0;
    assign fifo_intf_2189.finish = finish;
    csv_file_dump fifo_csv_dumper_2189;
    csv_file_dump cstatus_csv_dumper_2189;
    df_fifo_monitor fifo_monitor_2189;
    df_fifo_intf fifo_intf_2190(clock,reset);
    assign fifo_intf_2190.rd_en = AESL_inst_myproject.layer3_out_837_U.if_read & AESL_inst_myproject.layer3_out_837_U.if_empty_n;
    assign fifo_intf_2190.wr_en = AESL_inst_myproject.layer3_out_837_U.if_write & AESL_inst_myproject.layer3_out_837_U.if_full_n;
    assign fifo_intf_2190.fifo_rd_block = 0;
    assign fifo_intf_2190.fifo_wr_block = 0;
    assign fifo_intf_2190.finish = finish;
    csv_file_dump fifo_csv_dumper_2190;
    csv_file_dump cstatus_csv_dumper_2190;
    df_fifo_monitor fifo_monitor_2190;
    df_fifo_intf fifo_intf_2191(clock,reset);
    assign fifo_intf_2191.rd_en = AESL_inst_myproject.layer3_out_838_U.if_read & AESL_inst_myproject.layer3_out_838_U.if_empty_n;
    assign fifo_intf_2191.wr_en = AESL_inst_myproject.layer3_out_838_U.if_write & AESL_inst_myproject.layer3_out_838_U.if_full_n;
    assign fifo_intf_2191.fifo_rd_block = 0;
    assign fifo_intf_2191.fifo_wr_block = 0;
    assign fifo_intf_2191.finish = finish;
    csv_file_dump fifo_csv_dumper_2191;
    csv_file_dump cstatus_csv_dumper_2191;
    df_fifo_monitor fifo_monitor_2191;
    df_fifo_intf fifo_intf_2192(clock,reset);
    assign fifo_intf_2192.rd_en = AESL_inst_myproject.layer3_out_839_U.if_read & AESL_inst_myproject.layer3_out_839_U.if_empty_n;
    assign fifo_intf_2192.wr_en = AESL_inst_myproject.layer3_out_839_U.if_write & AESL_inst_myproject.layer3_out_839_U.if_full_n;
    assign fifo_intf_2192.fifo_rd_block = 0;
    assign fifo_intf_2192.fifo_wr_block = 0;
    assign fifo_intf_2192.finish = finish;
    csv_file_dump fifo_csv_dumper_2192;
    csv_file_dump cstatus_csv_dumper_2192;
    df_fifo_monitor fifo_monitor_2192;
    df_fifo_intf fifo_intf_2193(clock,reset);
    assign fifo_intf_2193.rd_en = AESL_inst_myproject.layer3_out_840_U.if_read & AESL_inst_myproject.layer3_out_840_U.if_empty_n;
    assign fifo_intf_2193.wr_en = AESL_inst_myproject.layer3_out_840_U.if_write & AESL_inst_myproject.layer3_out_840_U.if_full_n;
    assign fifo_intf_2193.fifo_rd_block = 0;
    assign fifo_intf_2193.fifo_wr_block = 0;
    assign fifo_intf_2193.finish = finish;
    csv_file_dump fifo_csv_dumper_2193;
    csv_file_dump cstatus_csv_dumper_2193;
    df_fifo_monitor fifo_monitor_2193;
    df_fifo_intf fifo_intf_2194(clock,reset);
    assign fifo_intf_2194.rd_en = AESL_inst_myproject.layer3_out_841_U.if_read & AESL_inst_myproject.layer3_out_841_U.if_empty_n;
    assign fifo_intf_2194.wr_en = AESL_inst_myproject.layer3_out_841_U.if_write & AESL_inst_myproject.layer3_out_841_U.if_full_n;
    assign fifo_intf_2194.fifo_rd_block = 0;
    assign fifo_intf_2194.fifo_wr_block = 0;
    assign fifo_intf_2194.finish = finish;
    csv_file_dump fifo_csv_dumper_2194;
    csv_file_dump cstatus_csv_dumper_2194;
    df_fifo_monitor fifo_monitor_2194;
    df_fifo_intf fifo_intf_2195(clock,reset);
    assign fifo_intf_2195.rd_en = AESL_inst_myproject.layer3_out_842_U.if_read & AESL_inst_myproject.layer3_out_842_U.if_empty_n;
    assign fifo_intf_2195.wr_en = AESL_inst_myproject.layer3_out_842_U.if_write & AESL_inst_myproject.layer3_out_842_U.if_full_n;
    assign fifo_intf_2195.fifo_rd_block = 0;
    assign fifo_intf_2195.fifo_wr_block = 0;
    assign fifo_intf_2195.finish = finish;
    csv_file_dump fifo_csv_dumper_2195;
    csv_file_dump cstatus_csv_dumper_2195;
    df_fifo_monitor fifo_monitor_2195;
    df_fifo_intf fifo_intf_2196(clock,reset);
    assign fifo_intf_2196.rd_en = AESL_inst_myproject.layer3_out_843_U.if_read & AESL_inst_myproject.layer3_out_843_U.if_empty_n;
    assign fifo_intf_2196.wr_en = AESL_inst_myproject.layer3_out_843_U.if_write & AESL_inst_myproject.layer3_out_843_U.if_full_n;
    assign fifo_intf_2196.fifo_rd_block = 0;
    assign fifo_intf_2196.fifo_wr_block = 0;
    assign fifo_intf_2196.finish = finish;
    csv_file_dump fifo_csv_dumper_2196;
    csv_file_dump cstatus_csv_dumper_2196;
    df_fifo_monitor fifo_monitor_2196;
    df_fifo_intf fifo_intf_2197(clock,reset);
    assign fifo_intf_2197.rd_en = AESL_inst_myproject.layer3_out_844_U.if_read & AESL_inst_myproject.layer3_out_844_U.if_empty_n;
    assign fifo_intf_2197.wr_en = AESL_inst_myproject.layer3_out_844_U.if_write & AESL_inst_myproject.layer3_out_844_U.if_full_n;
    assign fifo_intf_2197.fifo_rd_block = 0;
    assign fifo_intf_2197.fifo_wr_block = 0;
    assign fifo_intf_2197.finish = finish;
    csv_file_dump fifo_csv_dumper_2197;
    csv_file_dump cstatus_csv_dumper_2197;
    df_fifo_monitor fifo_monitor_2197;
    df_fifo_intf fifo_intf_2198(clock,reset);
    assign fifo_intf_2198.rd_en = AESL_inst_myproject.layer3_out_845_U.if_read & AESL_inst_myproject.layer3_out_845_U.if_empty_n;
    assign fifo_intf_2198.wr_en = AESL_inst_myproject.layer3_out_845_U.if_write & AESL_inst_myproject.layer3_out_845_U.if_full_n;
    assign fifo_intf_2198.fifo_rd_block = 0;
    assign fifo_intf_2198.fifo_wr_block = 0;
    assign fifo_intf_2198.finish = finish;
    csv_file_dump fifo_csv_dumper_2198;
    csv_file_dump cstatus_csv_dumper_2198;
    df_fifo_monitor fifo_monitor_2198;
    df_fifo_intf fifo_intf_2199(clock,reset);
    assign fifo_intf_2199.rd_en = AESL_inst_myproject.layer3_out_846_U.if_read & AESL_inst_myproject.layer3_out_846_U.if_empty_n;
    assign fifo_intf_2199.wr_en = AESL_inst_myproject.layer3_out_846_U.if_write & AESL_inst_myproject.layer3_out_846_U.if_full_n;
    assign fifo_intf_2199.fifo_rd_block = 0;
    assign fifo_intf_2199.fifo_wr_block = 0;
    assign fifo_intf_2199.finish = finish;
    csv_file_dump fifo_csv_dumper_2199;
    csv_file_dump cstatus_csv_dumper_2199;
    df_fifo_monitor fifo_monitor_2199;
    df_fifo_intf fifo_intf_2200(clock,reset);
    assign fifo_intf_2200.rd_en = AESL_inst_myproject.layer3_out_847_U.if_read & AESL_inst_myproject.layer3_out_847_U.if_empty_n;
    assign fifo_intf_2200.wr_en = AESL_inst_myproject.layer3_out_847_U.if_write & AESL_inst_myproject.layer3_out_847_U.if_full_n;
    assign fifo_intf_2200.fifo_rd_block = 0;
    assign fifo_intf_2200.fifo_wr_block = 0;
    assign fifo_intf_2200.finish = finish;
    csv_file_dump fifo_csv_dumper_2200;
    csv_file_dump cstatus_csv_dumper_2200;
    df_fifo_monitor fifo_monitor_2200;
    df_fifo_intf fifo_intf_2201(clock,reset);
    assign fifo_intf_2201.rd_en = AESL_inst_myproject.layer3_out_848_U.if_read & AESL_inst_myproject.layer3_out_848_U.if_empty_n;
    assign fifo_intf_2201.wr_en = AESL_inst_myproject.layer3_out_848_U.if_write & AESL_inst_myproject.layer3_out_848_U.if_full_n;
    assign fifo_intf_2201.fifo_rd_block = 0;
    assign fifo_intf_2201.fifo_wr_block = 0;
    assign fifo_intf_2201.finish = finish;
    csv_file_dump fifo_csv_dumper_2201;
    csv_file_dump cstatus_csv_dumper_2201;
    df_fifo_monitor fifo_monitor_2201;
    df_fifo_intf fifo_intf_2202(clock,reset);
    assign fifo_intf_2202.rd_en = AESL_inst_myproject.layer3_out_849_U.if_read & AESL_inst_myproject.layer3_out_849_U.if_empty_n;
    assign fifo_intf_2202.wr_en = AESL_inst_myproject.layer3_out_849_U.if_write & AESL_inst_myproject.layer3_out_849_U.if_full_n;
    assign fifo_intf_2202.fifo_rd_block = 0;
    assign fifo_intf_2202.fifo_wr_block = 0;
    assign fifo_intf_2202.finish = finish;
    csv_file_dump fifo_csv_dumper_2202;
    csv_file_dump cstatus_csv_dumper_2202;
    df_fifo_monitor fifo_monitor_2202;
    df_fifo_intf fifo_intf_2203(clock,reset);
    assign fifo_intf_2203.rd_en = AESL_inst_myproject.layer3_out_850_U.if_read & AESL_inst_myproject.layer3_out_850_U.if_empty_n;
    assign fifo_intf_2203.wr_en = AESL_inst_myproject.layer3_out_850_U.if_write & AESL_inst_myproject.layer3_out_850_U.if_full_n;
    assign fifo_intf_2203.fifo_rd_block = 0;
    assign fifo_intf_2203.fifo_wr_block = 0;
    assign fifo_intf_2203.finish = finish;
    csv_file_dump fifo_csv_dumper_2203;
    csv_file_dump cstatus_csv_dumper_2203;
    df_fifo_monitor fifo_monitor_2203;
    df_fifo_intf fifo_intf_2204(clock,reset);
    assign fifo_intf_2204.rd_en = AESL_inst_myproject.layer3_out_851_U.if_read & AESL_inst_myproject.layer3_out_851_U.if_empty_n;
    assign fifo_intf_2204.wr_en = AESL_inst_myproject.layer3_out_851_U.if_write & AESL_inst_myproject.layer3_out_851_U.if_full_n;
    assign fifo_intf_2204.fifo_rd_block = 0;
    assign fifo_intf_2204.fifo_wr_block = 0;
    assign fifo_intf_2204.finish = finish;
    csv_file_dump fifo_csv_dumper_2204;
    csv_file_dump cstatus_csv_dumper_2204;
    df_fifo_monitor fifo_monitor_2204;
    df_fifo_intf fifo_intf_2205(clock,reset);
    assign fifo_intf_2205.rd_en = AESL_inst_myproject.layer3_out_852_U.if_read & AESL_inst_myproject.layer3_out_852_U.if_empty_n;
    assign fifo_intf_2205.wr_en = AESL_inst_myproject.layer3_out_852_U.if_write & AESL_inst_myproject.layer3_out_852_U.if_full_n;
    assign fifo_intf_2205.fifo_rd_block = 0;
    assign fifo_intf_2205.fifo_wr_block = 0;
    assign fifo_intf_2205.finish = finish;
    csv_file_dump fifo_csv_dumper_2205;
    csv_file_dump cstatus_csv_dumper_2205;
    df_fifo_monitor fifo_monitor_2205;
    df_fifo_intf fifo_intf_2206(clock,reset);
    assign fifo_intf_2206.rd_en = AESL_inst_myproject.layer3_out_853_U.if_read & AESL_inst_myproject.layer3_out_853_U.if_empty_n;
    assign fifo_intf_2206.wr_en = AESL_inst_myproject.layer3_out_853_U.if_write & AESL_inst_myproject.layer3_out_853_U.if_full_n;
    assign fifo_intf_2206.fifo_rd_block = 0;
    assign fifo_intf_2206.fifo_wr_block = 0;
    assign fifo_intf_2206.finish = finish;
    csv_file_dump fifo_csv_dumper_2206;
    csv_file_dump cstatus_csv_dumper_2206;
    df_fifo_monitor fifo_monitor_2206;
    df_fifo_intf fifo_intf_2207(clock,reset);
    assign fifo_intf_2207.rd_en = AESL_inst_myproject.layer3_out_854_U.if_read & AESL_inst_myproject.layer3_out_854_U.if_empty_n;
    assign fifo_intf_2207.wr_en = AESL_inst_myproject.layer3_out_854_U.if_write & AESL_inst_myproject.layer3_out_854_U.if_full_n;
    assign fifo_intf_2207.fifo_rd_block = 0;
    assign fifo_intf_2207.fifo_wr_block = 0;
    assign fifo_intf_2207.finish = finish;
    csv_file_dump fifo_csv_dumper_2207;
    csv_file_dump cstatus_csv_dumper_2207;
    df_fifo_monitor fifo_monitor_2207;
    df_fifo_intf fifo_intf_2208(clock,reset);
    assign fifo_intf_2208.rd_en = AESL_inst_myproject.layer3_out_855_U.if_read & AESL_inst_myproject.layer3_out_855_U.if_empty_n;
    assign fifo_intf_2208.wr_en = AESL_inst_myproject.layer3_out_855_U.if_write & AESL_inst_myproject.layer3_out_855_U.if_full_n;
    assign fifo_intf_2208.fifo_rd_block = 0;
    assign fifo_intf_2208.fifo_wr_block = 0;
    assign fifo_intf_2208.finish = finish;
    csv_file_dump fifo_csv_dumper_2208;
    csv_file_dump cstatus_csv_dumper_2208;
    df_fifo_monitor fifo_monitor_2208;
    df_fifo_intf fifo_intf_2209(clock,reset);
    assign fifo_intf_2209.rd_en = AESL_inst_myproject.layer3_out_856_U.if_read & AESL_inst_myproject.layer3_out_856_U.if_empty_n;
    assign fifo_intf_2209.wr_en = AESL_inst_myproject.layer3_out_856_U.if_write & AESL_inst_myproject.layer3_out_856_U.if_full_n;
    assign fifo_intf_2209.fifo_rd_block = 0;
    assign fifo_intf_2209.fifo_wr_block = 0;
    assign fifo_intf_2209.finish = finish;
    csv_file_dump fifo_csv_dumper_2209;
    csv_file_dump cstatus_csv_dumper_2209;
    df_fifo_monitor fifo_monitor_2209;
    df_fifo_intf fifo_intf_2210(clock,reset);
    assign fifo_intf_2210.rd_en = AESL_inst_myproject.layer3_out_857_U.if_read & AESL_inst_myproject.layer3_out_857_U.if_empty_n;
    assign fifo_intf_2210.wr_en = AESL_inst_myproject.layer3_out_857_U.if_write & AESL_inst_myproject.layer3_out_857_U.if_full_n;
    assign fifo_intf_2210.fifo_rd_block = 0;
    assign fifo_intf_2210.fifo_wr_block = 0;
    assign fifo_intf_2210.finish = finish;
    csv_file_dump fifo_csv_dumper_2210;
    csv_file_dump cstatus_csv_dumper_2210;
    df_fifo_monitor fifo_monitor_2210;
    df_fifo_intf fifo_intf_2211(clock,reset);
    assign fifo_intf_2211.rd_en = AESL_inst_myproject.layer3_out_858_U.if_read & AESL_inst_myproject.layer3_out_858_U.if_empty_n;
    assign fifo_intf_2211.wr_en = AESL_inst_myproject.layer3_out_858_U.if_write & AESL_inst_myproject.layer3_out_858_U.if_full_n;
    assign fifo_intf_2211.fifo_rd_block = 0;
    assign fifo_intf_2211.fifo_wr_block = 0;
    assign fifo_intf_2211.finish = finish;
    csv_file_dump fifo_csv_dumper_2211;
    csv_file_dump cstatus_csv_dumper_2211;
    df_fifo_monitor fifo_monitor_2211;
    df_fifo_intf fifo_intf_2212(clock,reset);
    assign fifo_intf_2212.rd_en = AESL_inst_myproject.layer3_out_859_U.if_read & AESL_inst_myproject.layer3_out_859_U.if_empty_n;
    assign fifo_intf_2212.wr_en = AESL_inst_myproject.layer3_out_859_U.if_write & AESL_inst_myproject.layer3_out_859_U.if_full_n;
    assign fifo_intf_2212.fifo_rd_block = 0;
    assign fifo_intf_2212.fifo_wr_block = 0;
    assign fifo_intf_2212.finish = finish;
    csv_file_dump fifo_csv_dumper_2212;
    csv_file_dump cstatus_csv_dumper_2212;
    df_fifo_monitor fifo_monitor_2212;
    df_fifo_intf fifo_intf_2213(clock,reset);
    assign fifo_intf_2213.rd_en = AESL_inst_myproject.layer3_out_860_U.if_read & AESL_inst_myproject.layer3_out_860_U.if_empty_n;
    assign fifo_intf_2213.wr_en = AESL_inst_myproject.layer3_out_860_U.if_write & AESL_inst_myproject.layer3_out_860_U.if_full_n;
    assign fifo_intf_2213.fifo_rd_block = 0;
    assign fifo_intf_2213.fifo_wr_block = 0;
    assign fifo_intf_2213.finish = finish;
    csv_file_dump fifo_csv_dumper_2213;
    csv_file_dump cstatus_csv_dumper_2213;
    df_fifo_monitor fifo_monitor_2213;
    df_fifo_intf fifo_intf_2214(clock,reset);
    assign fifo_intf_2214.rd_en = AESL_inst_myproject.layer3_out_861_U.if_read & AESL_inst_myproject.layer3_out_861_U.if_empty_n;
    assign fifo_intf_2214.wr_en = AESL_inst_myproject.layer3_out_861_U.if_write & AESL_inst_myproject.layer3_out_861_U.if_full_n;
    assign fifo_intf_2214.fifo_rd_block = 0;
    assign fifo_intf_2214.fifo_wr_block = 0;
    assign fifo_intf_2214.finish = finish;
    csv_file_dump fifo_csv_dumper_2214;
    csv_file_dump cstatus_csv_dumper_2214;
    df_fifo_monitor fifo_monitor_2214;
    df_fifo_intf fifo_intf_2215(clock,reset);
    assign fifo_intf_2215.rd_en = AESL_inst_myproject.layer3_out_862_U.if_read & AESL_inst_myproject.layer3_out_862_U.if_empty_n;
    assign fifo_intf_2215.wr_en = AESL_inst_myproject.layer3_out_862_U.if_write & AESL_inst_myproject.layer3_out_862_U.if_full_n;
    assign fifo_intf_2215.fifo_rd_block = 0;
    assign fifo_intf_2215.fifo_wr_block = 0;
    assign fifo_intf_2215.finish = finish;
    csv_file_dump fifo_csv_dumper_2215;
    csv_file_dump cstatus_csv_dumper_2215;
    df_fifo_monitor fifo_monitor_2215;
    df_fifo_intf fifo_intf_2216(clock,reset);
    assign fifo_intf_2216.rd_en = AESL_inst_myproject.layer3_out_863_U.if_read & AESL_inst_myproject.layer3_out_863_U.if_empty_n;
    assign fifo_intf_2216.wr_en = AESL_inst_myproject.layer3_out_863_U.if_write & AESL_inst_myproject.layer3_out_863_U.if_full_n;
    assign fifo_intf_2216.fifo_rd_block = 0;
    assign fifo_intf_2216.fifo_wr_block = 0;
    assign fifo_intf_2216.finish = finish;
    csv_file_dump fifo_csv_dumper_2216;
    csv_file_dump cstatus_csv_dumper_2216;
    df_fifo_monitor fifo_monitor_2216;
    df_fifo_intf fifo_intf_2217(clock,reset);
    assign fifo_intf_2217.rd_en = AESL_inst_myproject.layer3_out_864_U.if_read & AESL_inst_myproject.layer3_out_864_U.if_empty_n;
    assign fifo_intf_2217.wr_en = AESL_inst_myproject.layer3_out_864_U.if_write & AESL_inst_myproject.layer3_out_864_U.if_full_n;
    assign fifo_intf_2217.fifo_rd_block = 0;
    assign fifo_intf_2217.fifo_wr_block = 0;
    assign fifo_intf_2217.finish = finish;
    csv_file_dump fifo_csv_dumper_2217;
    csv_file_dump cstatus_csv_dumper_2217;
    df_fifo_monitor fifo_monitor_2217;
    df_fifo_intf fifo_intf_2218(clock,reset);
    assign fifo_intf_2218.rd_en = AESL_inst_myproject.layer3_out_865_U.if_read & AESL_inst_myproject.layer3_out_865_U.if_empty_n;
    assign fifo_intf_2218.wr_en = AESL_inst_myproject.layer3_out_865_U.if_write & AESL_inst_myproject.layer3_out_865_U.if_full_n;
    assign fifo_intf_2218.fifo_rd_block = 0;
    assign fifo_intf_2218.fifo_wr_block = 0;
    assign fifo_intf_2218.finish = finish;
    csv_file_dump fifo_csv_dumper_2218;
    csv_file_dump cstatus_csv_dumper_2218;
    df_fifo_monitor fifo_monitor_2218;
    df_fifo_intf fifo_intf_2219(clock,reset);
    assign fifo_intf_2219.rd_en = AESL_inst_myproject.layer3_out_866_U.if_read & AESL_inst_myproject.layer3_out_866_U.if_empty_n;
    assign fifo_intf_2219.wr_en = AESL_inst_myproject.layer3_out_866_U.if_write & AESL_inst_myproject.layer3_out_866_U.if_full_n;
    assign fifo_intf_2219.fifo_rd_block = 0;
    assign fifo_intf_2219.fifo_wr_block = 0;
    assign fifo_intf_2219.finish = finish;
    csv_file_dump fifo_csv_dumper_2219;
    csv_file_dump cstatus_csv_dumper_2219;
    df_fifo_monitor fifo_monitor_2219;
    df_fifo_intf fifo_intf_2220(clock,reset);
    assign fifo_intf_2220.rd_en = AESL_inst_myproject.layer3_out_867_U.if_read & AESL_inst_myproject.layer3_out_867_U.if_empty_n;
    assign fifo_intf_2220.wr_en = AESL_inst_myproject.layer3_out_867_U.if_write & AESL_inst_myproject.layer3_out_867_U.if_full_n;
    assign fifo_intf_2220.fifo_rd_block = 0;
    assign fifo_intf_2220.fifo_wr_block = 0;
    assign fifo_intf_2220.finish = finish;
    csv_file_dump fifo_csv_dumper_2220;
    csv_file_dump cstatus_csv_dumper_2220;
    df_fifo_monitor fifo_monitor_2220;
    df_fifo_intf fifo_intf_2221(clock,reset);
    assign fifo_intf_2221.rd_en = AESL_inst_myproject.layer3_out_868_U.if_read & AESL_inst_myproject.layer3_out_868_U.if_empty_n;
    assign fifo_intf_2221.wr_en = AESL_inst_myproject.layer3_out_868_U.if_write & AESL_inst_myproject.layer3_out_868_U.if_full_n;
    assign fifo_intf_2221.fifo_rd_block = 0;
    assign fifo_intf_2221.fifo_wr_block = 0;
    assign fifo_intf_2221.finish = finish;
    csv_file_dump fifo_csv_dumper_2221;
    csv_file_dump cstatus_csv_dumper_2221;
    df_fifo_monitor fifo_monitor_2221;
    df_fifo_intf fifo_intf_2222(clock,reset);
    assign fifo_intf_2222.rd_en = AESL_inst_myproject.layer3_out_869_U.if_read & AESL_inst_myproject.layer3_out_869_U.if_empty_n;
    assign fifo_intf_2222.wr_en = AESL_inst_myproject.layer3_out_869_U.if_write & AESL_inst_myproject.layer3_out_869_U.if_full_n;
    assign fifo_intf_2222.fifo_rd_block = 0;
    assign fifo_intf_2222.fifo_wr_block = 0;
    assign fifo_intf_2222.finish = finish;
    csv_file_dump fifo_csv_dumper_2222;
    csv_file_dump cstatus_csv_dumper_2222;
    df_fifo_monitor fifo_monitor_2222;
    df_fifo_intf fifo_intf_2223(clock,reset);
    assign fifo_intf_2223.rd_en = AESL_inst_myproject.layer3_out_870_U.if_read & AESL_inst_myproject.layer3_out_870_U.if_empty_n;
    assign fifo_intf_2223.wr_en = AESL_inst_myproject.layer3_out_870_U.if_write & AESL_inst_myproject.layer3_out_870_U.if_full_n;
    assign fifo_intf_2223.fifo_rd_block = 0;
    assign fifo_intf_2223.fifo_wr_block = 0;
    assign fifo_intf_2223.finish = finish;
    csv_file_dump fifo_csv_dumper_2223;
    csv_file_dump cstatus_csv_dumper_2223;
    df_fifo_monitor fifo_monitor_2223;
    df_fifo_intf fifo_intf_2224(clock,reset);
    assign fifo_intf_2224.rd_en = AESL_inst_myproject.layer3_out_871_U.if_read & AESL_inst_myproject.layer3_out_871_U.if_empty_n;
    assign fifo_intf_2224.wr_en = AESL_inst_myproject.layer3_out_871_U.if_write & AESL_inst_myproject.layer3_out_871_U.if_full_n;
    assign fifo_intf_2224.fifo_rd_block = 0;
    assign fifo_intf_2224.fifo_wr_block = 0;
    assign fifo_intf_2224.finish = finish;
    csv_file_dump fifo_csv_dumper_2224;
    csv_file_dump cstatus_csv_dumper_2224;
    df_fifo_monitor fifo_monitor_2224;
    df_fifo_intf fifo_intf_2225(clock,reset);
    assign fifo_intf_2225.rd_en = AESL_inst_myproject.layer3_out_872_U.if_read & AESL_inst_myproject.layer3_out_872_U.if_empty_n;
    assign fifo_intf_2225.wr_en = AESL_inst_myproject.layer3_out_872_U.if_write & AESL_inst_myproject.layer3_out_872_U.if_full_n;
    assign fifo_intf_2225.fifo_rd_block = 0;
    assign fifo_intf_2225.fifo_wr_block = 0;
    assign fifo_intf_2225.finish = finish;
    csv_file_dump fifo_csv_dumper_2225;
    csv_file_dump cstatus_csv_dumper_2225;
    df_fifo_monitor fifo_monitor_2225;
    df_fifo_intf fifo_intf_2226(clock,reset);
    assign fifo_intf_2226.rd_en = AESL_inst_myproject.layer3_out_873_U.if_read & AESL_inst_myproject.layer3_out_873_U.if_empty_n;
    assign fifo_intf_2226.wr_en = AESL_inst_myproject.layer3_out_873_U.if_write & AESL_inst_myproject.layer3_out_873_U.if_full_n;
    assign fifo_intf_2226.fifo_rd_block = 0;
    assign fifo_intf_2226.fifo_wr_block = 0;
    assign fifo_intf_2226.finish = finish;
    csv_file_dump fifo_csv_dumper_2226;
    csv_file_dump cstatus_csv_dumper_2226;
    df_fifo_monitor fifo_monitor_2226;
    df_fifo_intf fifo_intf_2227(clock,reset);
    assign fifo_intf_2227.rd_en = AESL_inst_myproject.layer3_out_874_U.if_read & AESL_inst_myproject.layer3_out_874_U.if_empty_n;
    assign fifo_intf_2227.wr_en = AESL_inst_myproject.layer3_out_874_U.if_write & AESL_inst_myproject.layer3_out_874_U.if_full_n;
    assign fifo_intf_2227.fifo_rd_block = 0;
    assign fifo_intf_2227.fifo_wr_block = 0;
    assign fifo_intf_2227.finish = finish;
    csv_file_dump fifo_csv_dumper_2227;
    csv_file_dump cstatus_csv_dumper_2227;
    df_fifo_monitor fifo_monitor_2227;
    df_fifo_intf fifo_intf_2228(clock,reset);
    assign fifo_intf_2228.rd_en = AESL_inst_myproject.layer3_out_875_U.if_read & AESL_inst_myproject.layer3_out_875_U.if_empty_n;
    assign fifo_intf_2228.wr_en = AESL_inst_myproject.layer3_out_875_U.if_write & AESL_inst_myproject.layer3_out_875_U.if_full_n;
    assign fifo_intf_2228.fifo_rd_block = 0;
    assign fifo_intf_2228.fifo_wr_block = 0;
    assign fifo_intf_2228.finish = finish;
    csv_file_dump fifo_csv_dumper_2228;
    csv_file_dump cstatus_csv_dumper_2228;
    df_fifo_monitor fifo_monitor_2228;
    df_fifo_intf fifo_intf_2229(clock,reset);
    assign fifo_intf_2229.rd_en = AESL_inst_myproject.layer3_out_876_U.if_read & AESL_inst_myproject.layer3_out_876_U.if_empty_n;
    assign fifo_intf_2229.wr_en = AESL_inst_myproject.layer3_out_876_U.if_write & AESL_inst_myproject.layer3_out_876_U.if_full_n;
    assign fifo_intf_2229.fifo_rd_block = 0;
    assign fifo_intf_2229.fifo_wr_block = 0;
    assign fifo_intf_2229.finish = finish;
    csv_file_dump fifo_csv_dumper_2229;
    csv_file_dump cstatus_csv_dumper_2229;
    df_fifo_monitor fifo_monitor_2229;
    df_fifo_intf fifo_intf_2230(clock,reset);
    assign fifo_intf_2230.rd_en = AESL_inst_myproject.layer3_out_877_U.if_read & AESL_inst_myproject.layer3_out_877_U.if_empty_n;
    assign fifo_intf_2230.wr_en = AESL_inst_myproject.layer3_out_877_U.if_write & AESL_inst_myproject.layer3_out_877_U.if_full_n;
    assign fifo_intf_2230.fifo_rd_block = 0;
    assign fifo_intf_2230.fifo_wr_block = 0;
    assign fifo_intf_2230.finish = finish;
    csv_file_dump fifo_csv_dumper_2230;
    csv_file_dump cstatus_csv_dumper_2230;
    df_fifo_monitor fifo_monitor_2230;
    df_fifo_intf fifo_intf_2231(clock,reset);
    assign fifo_intf_2231.rd_en = AESL_inst_myproject.layer3_out_878_U.if_read & AESL_inst_myproject.layer3_out_878_U.if_empty_n;
    assign fifo_intf_2231.wr_en = AESL_inst_myproject.layer3_out_878_U.if_write & AESL_inst_myproject.layer3_out_878_U.if_full_n;
    assign fifo_intf_2231.fifo_rd_block = 0;
    assign fifo_intf_2231.fifo_wr_block = 0;
    assign fifo_intf_2231.finish = finish;
    csv_file_dump fifo_csv_dumper_2231;
    csv_file_dump cstatus_csv_dumper_2231;
    df_fifo_monitor fifo_monitor_2231;
    df_fifo_intf fifo_intf_2232(clock,reset);
    assign fifo_intf_2232.rd_en = AESL_inst_myproject.layer3_out_879_U.if_read & AESL_inst_myproject.layer3_out_879_U.if_empty_n;
    assign fifo_intf_2232.wr_en = AESL_inst_myproject.layer3_out_879_U.if_write & AESL_inst_myproject.layer3_out_879_U.if_full_n;
    assign fifo_intf_2232.fifo_rd_block = 0;
    assign fifo_intf_2232.fifo_wr_block = 0;
    assign fifo_intf_2232.finish = finish;
    csv_file_dump fifo_csv_dumper_2232;
    csv_file_dump cstatus_csv_dumper_2232;
    df_fifo_monitor fifo_monitor_2232;
    df_fifo_intf fifo_intf_2233(clock,reset);
    assign fifo_intf_2233.rd_en = AESL_inst_myproject.layer3_out_880_U.if_read & AESL_inst_myproject.layer3_out_880_U.if_empty_n;
    assign fifo_intf_2233.wr_en = AESL_inst_myproject.layer3_out_880_U.if_write & AESL_inst_myproject.layer3_out_880_U.if_full_n;
    assign fifo_intf_2233.fifo_rd_block = 0;
    assign fifo_intf_2233.fifo_wr_block = 0;
    assign fifo_intf_2233.finish = finish;
    csv_file_dump fifo_csv_dumper_2233;
    csv_file_dump cstatus_csv_dumper_2233;
    df_fifo_monitor fifo_monitor_2233;
    df_fifo_intf fifo_intf_2234(clock,reset);
    assign fifo_intf_2234.rd_en = AESL_inst_myproject.layer3_out_881_U.if_read & AESL_inst_myproject.layer3_out_881_U.if_empty_n;
    assign fifo_intf_2234.wr_en = AESL_inst_myproject.layer3_out_881_U.if_write & AESL_inst_myproject.layer3_out_881_U.if_full_n;
    assign fifo_intf_2234.fifo_rd_block = 0;
    assign fifo_intf_2234.fifo_wr_block = 0;
    assign fifo_intf_2234.finish = finish;
    csv_file_dump fifo_csv_dumper_2234;
    csv_file_dump cstatus_csv_dumper_2234;
    df_fifo_monitor fifo_monitor_2234;
    df_fifo_intf fifo_intf_2235(clock,reset);
    assign fifo_intf_2235.rd_en = AESL_inst_myproject.layer3_out_882_U.if_read & AESL_inst_myproject.layer3_out_882_U.if_empty_n;
    assign fifo_intf_2235.wr_en = AESL_inst_myproject.layer3_out_882_U.if_write & AESL_inst_myproject.layer3_out_882_U.if_full_n;
    assign fifo_intf_2235.fifo_rd_block = 0;
    assign fifo_intf_2235.fifo_wr_block = 0;
    assign fifo_intf_2235.finish = finish;
    csv_file_dump fifo_csv_dumper_2235;
    csv_file_dump cstatus_csv_dumper_2235;
    df_fifo_monitor fifo_monitor_2235;
    df_fifo_intf fifo_intf_2236(clock,reset);
    assign fifo_intf_2236.rd_en = AESL_inst_myproject.layer3_out_883_U.if_read & AESL_inst_myproject.layer3_out_883_U.if_empty_n;
    assign fifo_intf_2236.wr_en = AESL_inst_myproject.layer3_out_883_U.if_write & AESL_inst_myproject.layer3_out_883_U.if_full_n;
    assign fifo_intf_2236.fifo_rd_block = 0;
    assign fifo_intf_2236.fifo_wr_block = 0;
    assign fifo_intf_2236.finish = finish;
    csv_file_dump fifo_csv_dumper_2236;
    csv_file_dump cstatus_csv_dumper_2236;
    df_fifo_monitor fifo_monitor_2236;
    df_fifo_intf fifo_intf_2237(clock,reset);
    assign fifo_intf_2237.rd_en = AESL_inst_myproject.layer3_out_884_U.if_read & AESL_inst_myproject.layer3_out_884_U.if_empty_n;
    assign fifo_intf_2237.wr_en = AESL_inst_myproject.layer3_out_884_U.if_write & AESL_inst_myproject.layer3_out_884_U.if_full_n;
    assign fifo_intf_2237.fifo_rd_block = 0;
    assign fifo_intf_2237.fifo_wr_block = 0;
    assign fifo_intf_2237.finish = finish;
    csv_file_dump fifo_csv_dumper_2237;
    csv_file_dump cstatus_csv_dumper_2237;
    df_fifo_monitor fifo_monitor_2237;
    df_fifo_intf fifo_intf_2238(clock,reset);
    assign fifo_intf_2238.rd_en = AESL_inst_myproject.layer3_out_885_U.if_read & AESL_inst_myproject.layer3_out_885_U.if_empty_n;
    assign fifo_intf_2238.wr_en = AESL_inst_myproject.layer3_out_885_U.if_write & AESL_inst_myproject.layer3_out_885_U.if_full_n;
    assign fifo_intf_2238.fifo_rd_block = 0;
    assign fifo_intf_2238.fifo_wr_block = 0;
    assign fifo_intf_2238.finish = finish;
    csv_file_dump fifo_csv_dumper_2238;
    csv_file_dump cstatus_csv_dumper_2238;
    df_fifo_monitor fifo_monitor_2238;
    df_fifo_intf fifo_intf_2239(clock,reset);
    assign fifo_intf_2239.rd_en = AESL_inst_myproject.layer3_out_886_U.if_read & AESL_inst_myproject.layer3_out_886_U.if_empty_n;
    assign fifo_intf_2239.wr_en = AESL_inst_myproject.layer3_out_886_U.if_write & AESL_inst_myproject.layer3_out_886_U.if_full_n;
    assign fifo_intf_2239.fifo_rd_block = 0;
    assign fifo_intf_2239.fifo_wr_block = 0;
    assign fifo_intf_2239.finish = finish;
    csv_file_dump fifo_csv_dumper_2239;
    csv_file_dump cstatus_csv_dumper_2239;
    df_fifo_monitor fifo_monitor_2239;
    df_fifo_intf fifo_intf_2240(clock,reset);
    assign fifo_intf_2240.rd_en = AESL_inst_myproject.layer3_out_887_U.if_read & AESL_inst_myproject.layer3_out_887_U.if_empty_n;
    assign fifo_intf_2240.wr_en = AESL_inst_myproject.layer3_out_887_U.if_write & AESL_inst_myproject.layer3_out_887_U.if_full_n;
    assign fifo_intf_2240.fifo_rd_block = 0;
    assign fifo_intf_2240.fifo_wr_block = 0;
    assign fifo_intf_2240.finish = finish;
    csv_file_dump fifo_csv_dumper_2240;
    csv_file_dump cstatus_csv_dumper_2240;
    df_fifo_monitor fifo_monitor_2240;
    df_fifo_intf fifo_intf_2241(clock,reset);
    assign fifo_intf_2241.rd_en = AESL_inst_myproject.layer3_out_888_U.if_read & AESL_inst_myproject.layer3_out_888_U.if_empty_n;
    assign fifo_intf_2241.wr_en = AESL_inst_myproject.layer3_out_888_U.if_write & AESL_inst_myproject.layer3_out_888_U.if_full_n;
    assign fifo_intf_2241.fifo_rd_block = 0;
    assign fifo_intf_2241.fifo_wr_block = 0;
    assign fifo_intf_2241.finish = finish;
    csv_file_dump fifo_csv_dumper_2241;
    csv_file_dump cstatus_csv_dumper_2241;
    df_fifo_monitor fifo_monitor_2241;
    df_fifo_intf fifo_intf_2242(clock,reset);
    assign fifo_intf_2242.rd_en = AESL_inst_myproject.layer3_out_889_U.if_read & AESL_inst_myproject.layer3_out_889_U.if_empty_n;
    assign fifo_intf_2242.wr_en = AESL_inst_myproject.layer3_out_889_U.if_write & AESL_inst_myproject.layer3_out_889_U.if_full_n;
    assign fifo_intf_2242.fifo_rd_block = 0;
    assign fifo_intf_2242.fifo_wr_block = 0;
    assign fifo_intf_2242.finish = finish;
    csv_file_dump fifo_csv_dumper_2242;
    csv_file_dump cstatus_csv_dumper_2242;
    df_fifo_monitor fifo_monitor_2242;
    df_fifo_intf fifo_intf_2243(clock,reset);
    assign fifo_intf_2243.rd_en = AESL_inst_myproject.layer3_out_890_U.if_read & AESL_inst_myproject.layer3_out_890_U.if_empty_n;
    assign fifo_intf_2243.wr_en = AESL_inst_myproject.layer3_out_890_U.if_write & AESL_inst_myproject.layer3_out_890_U.if_full_n;
    assign fifo_intf_2243.fifo_rd_block = 0;
    assign fifo_intf_2243.fifo_wr_block = 0;
    assign fifo_intf_2243.finish = finish;
    csv_file_dump fifo_csv_dumper_2243;
    csv_file_dump cstatus_csv_dumper_2243;
    df_fifo_monitor fifo_monitor_2243;
    df_fifo_intf fifo_intf_2244(clock,reset);
    assign fifo_intf_2244.rd_en = AESL_inst_myproject.layer3_out_891_U.if_read & AESL_inst_myproject.layer3_out_891_U.if_empty_n;
    assign fifo_intf_2244.wr_en = AESL_inst_myproject.layer3_out_891_U.if_write & AESL_inst_myproject.layer3_out_891_U.if_full_n;
    assign fifo_intf_2244.fifo_rd_block = 0;
    assign fifo_intf_2244.fifo_wr_block = 0;
    assign fifo_intf_2244.finish = finish;
    csv_file_dump fifo_csv_dumper_2244;
    csv_file_dump cstatus_csv_dumper_2244;
    df_fifo_monitor fifo_monitor_2244;
    df_fifo_intf fifo_intf_2245(clock,reset);
    assign fifo_intf_2245.rd_en = AESL_inst_myproject.layer3_out_892_U.if_read & AESL_inst_myproject.layer3_out_892_U.if_empty_n;
    assign fifo_intf_2245.wr_en = AESL_inst_myproject.layer3_out_892_U.if_write & AESL_inst_myproject.layer3_out_892_U.if_full_n;
    assign fifo_intf_2245.fifo_rd_block = 0;
    assign fifo_intf_2245.fifo_wr_block = 0;
    assign fifo_intf_2245.finish = finish;
    csv_file_dump fifo_csv_dumper_2245;
    csv_file_dump cstatus_csv_dumper_2245;
    df_fifo_monitor fifo_monitor_2245;
    df_fifo_intf fifo_intf_2246(clock,reset);
    assign fifo_intf_2246.rd_en = AESL_inst_myproject.layer3_out_893_U.if_read & AESL_inst_myproject.layer3_out_893_U.if_empty_n;
    assign fifo_intf_2246.wr_en = AESL_inst_myproject.layer3_out_893_U.if_write & AESL_inst_myproject.layer3_out_893_U.if_full_n;
    assign fifo_intf_2246.fifo_rd_block = 0;
    assign fifo_intf_2246.fifo_wr_block = 0;
    assign fifo_intf_2246.finish = finish;
    csv_file_dump fifo_csv_dumper_2246;
    csv_file_dump cstatus_csv_dumper_2246;
    df_fifo_monitor fifo_monitor_2246;
    df_fifo_intf fifo_intf_2247(clock,reset);
    assign fifo_intf_2247.rd_en = AESL_inst_myproject.layer3_out_894_U.if_read & AESL_inst_myproject.layer3_out_894_U.if_empty_n;
    assign fifo_intf_2247.wr_en = AESL_inst_myproject.layer3_out_894_U.if_write & AESL_inst_myproject.layer3_out_894_U.if_full_n;
    assign fifo_intf_2247.fifo_rd_block = 0;
    assign fifo_intf_2247.fifo_wr_block = 0;
    assign fifo_intf_2247.finish = finish;
    csv_file_dump fifo_csv_dumper_2247;
    csv_file_dump cstatus_csv_dumper_2247;
    df_fifo_monitor fifo_monitor_2247;
    df_fifo_intf fifo_intf_2248(clock,reset);
    assign fifo_intf_2248.rd_en = AESL_inst_myproject.layer3_out_895_U.if_read & AESL_inst_myproject.layer3_out_895_U.if_empty_n;
    assign fifo_intf_2248.wr_en = AESL_inst_myproject.layer3_out_895_U.if_write & AESL_inst_myproject.layer3_out_895_U.if_full_n;
    assign fifo_intf_2248.fifo_rd_block = 0;
    assign fifo_intf_2248.fifo_wr_block = 0;
    assign fifo_intf_2248.finish = finish;
    csv_file_dump fifo_csv_dumper_2248;
    csv_file_dump cstatus_csv_dumper_2248;
    df_fifo_monitor fifo_monitor_2248;
    df_fifo_intf fifo_intf_2249(clock,reset);
    assign fifo_intf_2249.rd_en = AESL_inst_myproject.layer3_out_896_U.if_read & AESL_inst_myproject.layer3_out_896_U.if_empty_n;
    assign fifo_intf_2249.wr_en = AESL_inst_myproject.layer3_out_896_U.if_write & AESL_inst_myproject.layer3_out_896_U.if_full_n;
    assign fifo_intf_2249.fifo_rd_block = 0;
    assign fifo_intf_2249.fifo_wr_block = 0;
    assign fifo_intf_2249.finish = finish;
    csv_file_dump fifo_csv_dumper_2249;
    csv_file_dump cstatus_csv_dumper_2249;
    df_fifo_monitor fifo_monitor_2249;
    df_fifo_intf fifo_intf_2250(clock,reset);
    assign fifo_intf_2250.rd_en = AESL_inst_myproject.layer3_out_897_U.if_read & AESL_inst_myproject.layer3_out_897_U.if_empty_n;
    assign fifo_intf_2250.wr_en = AESL_inst_myproject.layer3_out_897_U.if_write & AESL_inst_myproject.layer3_out_897_U.if_full_n;
    assign fifo_intf_2250.fifo_rd_block = 0;
    assign fifo_intf_2250.fifo_wr_block = 0;
    assign fifo_intf_2250.finish = finish;
    csv_file_dump fifo_csv_dumper_2250;
    csv_file_dump cstatus_csv_dumper_2250;
    df_fifo_monitor fifo_monitor_2250;
    df_fifo_intf fifo_intf_2251(clock,reset);
    assign fifo_intf_2251.rd_en = AESL_inst_myproject.layer3_out_898_U.if_read & AESL_inst_myproject.layer3_out_898_U.if_empty_n;
    assign fifo_intf_2251.wr_en = AESL_inst_myproject.layer3_out_898_U.if_write & AESL_inst_myproject.layer3_out_898_U.if_full_n;
    assign fifo_intf_2251.fifo_rd_block = 0;
    assign fifo_intf_2251.fifo_wr_block = 0;
    assign fifo_intf_2251.finish = finish;
    csv_file_dump fifo_csv_dumper_2251;
    csv_file_dump cstatus_csv_dumper_2251;
    df_fifo_monitor fifo_monitor_2251;
    df_fifo_intf fifo_intf_2252(clock,reset);
    assign fifo_intf_2252.rd_en = AESL_inst_myproject.layer3_out_899_U.if_read & AESL_inst_myproject.layer3_out_899_U.if_empty_n;
    assign fifo_intf_2252.wr_en = AESL_inst_myproject.layer3_out_899_U.if_write & AESL_inst_myproject.layer3_out_899_U.if_full_n;
    assign fifo_intf_2252.fifo_rd_block = 0;
    assign fifo_intf_2252.fifo_wr_block = 0;
    assign fifo_intf_2252.finish = finish;
    csv_file_dump fifo_csv_dumper_2252;
    csv_file_dump cstatus_csv_dumper_2252;
    df_fifo_monitor fifo_monitor_2252;
    df_fifo_intf fifo_intf_2253(clock,reset);
    assign fifo_intf_2253.rd_en = AESL_inst_myproject.layer3_out_900_U.if_read & AESL_inst_myproject.layer3_out_900_U.if_empty_n;
    assign fifo_intf_2253.wr_en = AESL_inst_myproject.layer3_out_900_U.if_write & AESL_inst_myproject.layer3_out_900_U.if_full_n;
    assign fifo_intf_2253.fifo_rd_block = 0;
    assign fifo_intf_2253.fifo_wr_block = 0;
    assign fifo_intf_2253.finish = finish;
    csv_file_dump fifo_csv_dumper_2253;
    csv_file_dump cstatus_csv_dumper_2253;
    df_fifo_monitor fifo_monitor_2253;
    df_fifo_intf fifo_intf_2254(clock,reset);
    assign fifo_intf_2254.rd_en = AESL_inst_myproject.layer3_out_901_U.if_read & AESL_inst_myproject.layer3_out_901_U.if_empty_n;
    assign fifo_intf_2254.wr_en = AESL_inst_myproject.layer3_out_901_U.if_write & AESL_inst_myproject.layer3_out_901_U.if_full_n;
    assign fifo_intf_2254.fifo_rd_block = 0;
    assign fifo_intf_2254.fifo_wr_block = 0;
    assign fifo_intf_2254.finish = finish;
    csv_file_dump fifo_csv_dumper_2254;
    csv_file_dump cstatus_csv_dumper_2254;
    df_fifo_monitor fifo_monitor_2254;
    df_fifo_intf fifo_intf_2255(clock,reset);
    assign fifo_intf_2255.rd_en = AESL_inst_myproject.layer3_out_902_U.if_read & AESL_inst_myproject.layer3_out_902_U.if_empty_n;
    assign fifo_intf_2255.wr_en = AESL_inst_myproject.layer3_out_902_U.if_write & AESL_inst_myproject.layer3_out_902_U.if_full_n;
    assign fifo_intf_2255.fifo_rd_block = 0;
    assign fifo_intf_2255.fifo_wr_block = 0;
    assign fifo_intf_2255.finish = finish;
    csv_file_dump fifo_csv_dumper_2255;
    csv_file_dump cstatus_csv_dumper_2255;
    df_fifo_monitor fifo_monitor_2255;
    df_fifo_intf fifo_intf_2256(clock,reset);
    assign fifo_intf_2256.rd_en = AESL_inst_myproject.layer3_out_903_U.if_read & AESL_inst_myproject.layer3_out_903_U.if_empty_n;
    assign fifo_intf_2256.wr_en = AESL_inst_myproject.layer3_out_903_U.if_write & AESL_inst_myproject.layer3_out_903_U.if_full_n;
    assign fifo_intf_2256.fifo_rd_block = 0;
    assign fifo_intf_2256.fifo_wr_block = 0;
    assign fifo_intf_2256.finish = finish;
    csv_file_dump fifo_csv_dumper_2256;
    csv_file_dump cstatus_csv_dumper_2256;
    df_fifo_monitor fifo_monitor_2256;
    df_fifo_intf fifo_intf_2257(clock,reset);
    assign fifo_intf_2257.rd_en = AESL_inst_myproject.layer3_out_904_U.if_read & AESL_inst_myproject.layer3_out_904_U.if_empty_n;
    assign fifo_intf_2257.wr_en = AESL_inst_myproject.layer3_out_904_U.if_write & AESL_inst_myproject.layer3_out_904_U.if_full_n;
    assign fifo_intf_2257.fifo_rd_block = 0;
    assign fifo_intf_2257.fifo_wr_block = 0;
    assign fifo_intf_2257.finish = finish;
    csv_file_dump fifo_csv_dumper_2257;
    csv_file_dump cstatus_csv_dumper_2257;
    df_fifo_monitor fifo_monitor_2257;
    df_fifo_intf fifo_intf_2258(clock,reset);
    assign fifo_intf_2258.rd_en = AESL_inst_myproject.layer3_out_905_U.if_read & AESL_inst_myproject.layer3_out_905_U.if_empty_n;
    assign fifo_intf_2258.wr_en = AESL_inst_myproject.layer3_out_905_U.if_write & AESL_inst_myproject.layer3_out_905_U.if_full_n;
    assign fifo_intf_2258.fifo_rd_block = 0;
    assign fifo_intf_2258.fifo_wr_block = 0;
    assign fifo_intf_2258.finish = finish;
    csv_file_dump fifo_csv_dumper_2258;
    csv_file_dump cstatus_csv_dumper_2258;
    df_fifo_monitor fifo_monitor_2258;
    df_fifo_intf fifo_intf_2259(clock,reset);
    assign fifo_intf_2259.rd_en = AESL_inst_myproject.layer3_out_906_U.if_read & AESL_inst_myproject.layer3_out_906_U.if_empty_n;
    assign fifo_intf_2259.wr_en = AESL_inst_myproject.layer3_out_906_U.if_write & AESL_inst_myproject.layer3_out_906_U.if_full_n;
    assign fifo_intf_2259.fifo_rd_block = 0;
    assign fifo_intf_2259.fifo_wr_block = 0;
    assign fifo_intf_2259.finish = finish;
    csv_file_dump fifo_csv_dumper_2259;
    csv_file_dump cstatus_csv_dumper_2259;
    df_fifo_monitor fifo_monitor_2259;
    df_fifo_intf fifo_intf_2260(clock,reset);
    assign fifo_intf_2260.rd_en = AESL_inst_myproject.layer3_out_907_U.if_read & AESL_inst_myproject.layer3_out_907_U.if_empty_n;
    assign fifo_intf_2260.wr_en = AESL_inst_myproject.layer3_out_907_U.if_write & AESL_inst_myproject.layer3_out_907_U.if_full_n;
    assign fifo_intf_2260.fifo_rd_block = 0;
    assign fifo_intf_2260.fifo_wr_block = 0;
    assign fifo_intf_2260.finish = finish;
    csv_file_dump fifo_csv_dumper_2260;
    csv_file_dump cstatus_csv_dumper_2260;
    df_fifo_monitor fifo_monitor_2260;
    df_fifo_intf fifo_intf_2261(clock,reset);
    assign fifo_intf_2261.rd_en = AESL_inst_myproject.layer3_out_908_U.if_read & AESL_inst_myproject.layer3_out_908_U.if_empty_n;
    assign fifo_intf_2261.wr_en = AESL_inst_myproject.layer3_out_908_U.if_write & AESL_inst_myproject.layer3_out_908_U.if_full_n;
    assign fifo_intf_2261.fifo_rd_block = 0;
    assign fifo_intf_2261.fifo_wr_block = 0;
    assign fifo_intf_2261.finish = finish;
    csv_file_dump fifo_csv_dumper_2261;
    csv_file_dump cstatus_csv_dumper_2261;
    df_fifo_monitor fifo_monitor_2261;
    df_fifo_intf fifo_intf_2262(clock,reset);
    assign fifo_intf_2262.rd_en = AESL_inst_myproject.layer3_out_909_U.if_read & AESL_inst_myproject.layer3_out_909_U.if_empty_n;
    assign fifo_intf_2262.wr_en = AESL_inst_myproject.layer3_out_909_U.if_write & AESL_inst_myproject.layer3_out_909_U.if_full_n;
    assign fifo_intf_2262.fifo_rd_block = 0;
    assign fifo_intf_2262.fifo_wr_block = 0;
    assign fifo_intf_2262.finish = finish;
    csv_file_dump fifo_csv_dumper_2262;
    csv_file_dump cstatus_csv_dumper_2262;
    df_fifo_monitor fifo_monitor_2262;
    df_fifo_intf fifo_intf_2263(clock,reset);
    assign fifo_intf_2263.rd_en = AESL_inst_myproject.layer3_out_910_U.if_read & AESL_inst_myproject.layer3_out_910_U.if_empty_n;
    assign fifo_intf_2263.wr_en = AESL_inst_myproject.layer3_out_910_U.if_write & AESL_inst_myproject.layer3_out_910_U.if_full_n;
    assign fifo_intf_2263.fifo_rd_block = 0;
    assign fifo_intf_2263.fifo_wr_block = 0;
    assign fifo_intf_2263.finish = finish;
    csv_file_dump fifo_csv_dumper_2263;
    csv_file_dump cstatus_csv_dumper_2263;
    df_fifo_monitor fifo_monitor_2263;
    df_fifo_intf fifo_intf_2264(clock,reset);
    assign fifo_intf_2264.rd_en = AESL_inst_myproject.layer3_out_911_U.if_read & AESL_inst_myproject.layer3_out_911_U.if_empty_n;
    assign fifo_intf_2264.wr_en = AESL_inst_myproject.layer3_out_911_U.if_write & AESL_inst_myproject.layer3_out_911_U.if_full_n;
    assign fifo_intf_2264.fifo_rd_block = 0;
    assign fifo_intf_2264.fifo_wr_block = 0;
    assign fifo_intf_2264.finish = finish;
    csv_file_dump fifo_csv_dumper_2264;
    csv_file_dump cstatus_csv_dumper_2264;
    df_fifo_monitor fifo_monitor_2264;
    df_fifo_intf fifo_intf_2265(clock,reset);
    assign fifo_intf_2265.rd_en = AESL_inst_myproject.layer3_out_912_U.if_read & AESL_inst_myproject.layer3_out_912_U.if_empty_n;
    assign fifo_intf_2265.wr_en = AESL_inst_myproject.layer3_out_912_U.if_write & AESL_inst_myproject.layer3_out_912_U.if_full_n;
    assign fifo_intf_2265.fifo_rd_block = 0;
    assign fifo_intf_2265.fifo_wr_block = 0;
    assign fifo_intf_2265.finish = finish;
    csv_file_dump fifo_csv_dumper_2265;
    csv_file_dump cstatus_csv_dumper_2265;
    df_fifo_monitor fifo_monitor_2265;
    df_fifo_intf fifo_intf_2266(clock,reset);
    assign fifo_intf_2266.rd_en = AESL_inst_myproject.layer3_out_913_U.if_read & AESL_inst_myproject.layer3_out_913_U.if_empty_n;
    assign fifo_intf_2266.wr_en = AESL_inst_myproject.layer3_out_913_U.if_write & AESL_inst_myproject.layer3_out_913_U.if_full_n;
    assign fifo_intf_2266.fifo_rd_block = 0;
    assign fifo_intf_2266.fifo_wr_block = 0;
    assign fifo_intf_2266.finish = finish;
    csv_file_dump fifo_csv_dumper_2266;
    csv_file_dump cstatus_csv_dumper_2266;
    df_fifo_monitor fifo_monitor_2266;
    df_fifo_intf fifo_intf_2267(clock,reset);
    assign fifo_intf_2267.rd_en = AESL_inst_myproject.layer3_out_914_U.if_read & AESL_inst_myproject.layer3_out_914_U.if_empty_n;
    assign fifo_intf_2267.wr_en = AESL_inst_myproject.layer3_out_914_U.if_write & AESL_inst_myproject.layer3_out_914_U.if_full_n;
    assign fifo_intf_2267.fifo_rd_block = 0;
    assign fifo_intf_2267.fifo_wr_block = 0;
    assign fifo_intf_2267.finish = finish;
    csv_file_dump fifo_csv_dumper_2267;
    csv_file_dump cstatus_csv_dumper_2267;
    df_fifo_monitor fifo_monitor_2267;
    df_fifo_intf fifo_intf_2268(clock,reset);
    assign fifo_intf_2268.rd_en = AESL_inst_myproject.layer3_out_915_U.if_read & AESL_inst_myproject.layer3_out_915_U.if_empty_n;
    assign fifo_intf_2268.wr_en = AESL_inst_myproject.layer3_out_915_U.if_write & AESL_inst_myproject.layer3_out_915_U.if_full_n;
    assign fifo_intf_2268.fifo_rd_block = 0;
    assign fifo_intf_2268.fifo_wr_block = 0;
    assign fifo_intf_2268.finish = finish;
    csv_file_dump fifo_csv_dumper_2268;
    csv_file_dump cstatus_csv_dumper_2268;
    df_fifo_monitor fifo_monitor_2268;
    df_fifo_intf fifo_intf_2269(clock,reset);
    assign fifo_intf_2269.rd_en = AESL_inst_myproject.layer3_out_916_U.if_read & AESL_inst_myproject.layer3_out_916_U.if_empty_n;
    assign fifo_intf_2269.wr_en = AESL_inst_myproject.layer3_out_916_U.if_write & AESL_inst_myproject.layer3_out_916_U.if_full_n;
    assign fifo_intf_2269.fifo_rd_block = 0;
    assign fifo_intf_2269.fifo_wr_block = 0;
    assign fifo_intf_2269.finish = finish;
    csv_file_dump fifo_csv_dumper_2269;
    csv_file_dump cstatus_csv_dumper_2269;
    df_fifo_monitor fifo_monitor_2269;
    df_fifo_intf fifo_intf_2270(clock,reset);
    assign fifo_intf_2270.rd_en = AESL_inst_myproject.layer3_out_917_U.if_read & AESL_inst_myproject.layer3_out_917_U.if_empty_n;
    assign fifo_intf_2270.wr_en = AESL_inst_myproject.layer3_out_917_U.if_write & AESL_inst_myproject.layer3_out_917_U.if_full_n;
    assign fifo_intf_2270.fifo_rd_block = 0;
    assign fifo_intf_2270.fifo_wr_block = 0;
    assign fifo_intf_2270.finish = finish;
    csv_file_dump fifo_csv_dumper_2270;
    csv_file_dump cstatus_csv_dumper_2270;
    df_fifo_monitor fifo_monitor_2270;
    df_fifo_intf fifo_intf_2271(clock,reset);
    assign fifo_intf_2271.rd_en = AESL_inst_myproject.layer3_out_918_U.if_read & AESL_inst_myproject.layer3_out_918_U.if_empty_n;
    assign fifo_intf_2271.wr_en = AESL_inst_myproject.layer3_out_918_U.if_write & AESL_inst_myproject.layer3_out_918_U.if_full_n;
    assign fifo_intf_2271.fifo_rd_block = 0;
    assign fifo_intf_2271.fifo_wr_block = 0;
    assign fifo_intf_2271.finish = finish;
    csv_file_dump fifo_csv_dumper_2271;
    csv_file_dump cstatus_csv_dumper_2271;
    df_fifo_monitor fifo_monitor_2271;
    df_fifo_intf fifo_intf_2272(clock,reset);
    assign fifo_intf_2272.rd_en = AESL_inst_myproject.layer3_out_919_U.if_read & AESL_inst_myproject.layer3_out_919_U.if_empty_n;
    assign fifo_intf_2272.wr_en = AESL_inst_myproject.layer3_out_919_U.if_write & AESL_inst_myproject.layer3_out_919_U.if_full_n;
    assign fifo_intf_2272.fifo_rd_block = 0;
    assign fifo_intf_2272.fifo_wr_block = 0;
    assign fifo_intf_2272.finish = finish;
    csv_file_dump fifo_csv_dumper_2272;
    csv_file_dump cstatus_csv_dumper_2272;
    df_fifo_monitor fifo_monitor_2272;
    df_fifo_intf fifo_intf_2273(clock,reset);
    assign fifo_intf_2273.rd_en = AESL_inst_myproject.layer3_out_920_U.if_read & AESL_inst_myproject.layer3_out_920_U.if_empty_n;
    assign fifo_intf_2273.wr_en = AESL_inst_myproject.layer3_out_920_U.if_write & AESL_inst_myproject.layer3_out_920_U.if_full_n;
    assign fifo_intf_2273.fifo_rd_block = 0;
    assign fifo_intf_2273.fifo_wr_block = 0;
    assign fifo_intf_2273.finish = finish;
    csv_file_dump fifo_csv_dumper_2273;
    csv_file_dump cstatus_csv_dumper_2273;
    df_fifo_monitor fifo_monitor_2273;
    df_fifo_intf fifo_intf_2274(clock,reset);
    assign fifo_intf_2274.rd_en = AESL_inst_myproject.layer3_out_921_U.if_read & AESL_inst_myproject.layer3_out_921_U.if_empty_n;
    assign fifo_intf_2274.wr_en = AESL_inst_myproject.layer3_out_921_U.if_write & AESL_inst_myproject.layer3_out_921_U.if_full_n;
    assign fifo_intf_2274.fifo_rd_block = 0;
    assign fifo_intf_2274.fifo_wr_block = 0;
    assign fifo_intf_2274.finish = finish;
    csv_file_dump fifo_csv_dumper_2274;
    csv_file_dump cstatus_csv_dumper_2274;
    df_fifo_monitor fifo_monitor_2274;
    df_fifo_intf fifo_intf_2275(clock,reset);
    assign fifo_intf_2275.rd_en = AESL_inst_myproject.layer3_out_922_U.if_read & AESL_inst_myproject.layer3_out_922_U.if_empty_n;
    assign fifo_intf_2275.wr_en = AESL_inst_myproject.layer3_out_922_U.if_write & AESL_inst_myproject.layer3_out_922_U.if_full_n;
    assign fifo_intf_2275.fifo_rd_block = 0;
    assign fifo_intf_2275.fifo_wr_block = 0;
    assign fifo_intf_2275.finish = finish;
    csv_file_dump fifo_csv_dumper_2275;
    csv_file_dump cstatus_csv_dumper_2275;
    df_fifo_monitor fifo_monitor_2275;
    df_fifo_intf fifo_intf_2276(clock,reset);
    assign fifo_intf_2276.rd_en = AESL_inst_myproject.layer3_out_923_U.if_read & AESL_inst_myproject.layer3_out_923_U.if_empty_n;
    assign fifo_intf_2276.wr_en = AESL_inst_myproject.layer3_out_923_U.if_write & AESL_inst_myproject.layer3_out_923_U.if_full_n;
    assign fifo_intf_2276.fifo_rd_block = 0;
    assign fifo_intf_2276.fifo_wr_block = 0;
    assign fifo_intf_2276.finish = finish;
    csv_file_dump fifo_csv_dumper_2276;
    csv_file_dump cstatus_csv_dumper_2276;
    df_fifo_monitor fifo_monitor_2276;
    df_fifo_intf fifo_intf_2277(clock,reset);
    assign fifo_intf_2277.rd_en = AESL_inst_myproject.layer3_out_924_U.if_read & AESL_inst_myproject.layer3_out_924_U.if_empty_n;
    assign fifo_intf_2277.wr_en = AESL_inst_myproject.layer3_out_924_U.if_write & AESL_inst_myproject.layer3_out_924_U.if_full_n;
    assign fifo_intf_2277.fifo_rd_block = 0;
    assign fifo_intf_2277.fifo_wr_block = 0;
    assign fifo_intf_2277.finish = finish;
    csv_file_dump fifo_csv_dumper_2277;
    csv_file_dump cstatus_csv_dumper_2277;
    df_fifo_monitor fifo_monitor_2277;
    df_fifo_intf fifo_intf_2278(clock,reset);
    assign fifo_intf_2278.rd_en = AESL_inst_myproject.layer3_out_925_U.if_read & AESL_inst_myproject.layer3_out_925_U.if_empty_n;
    assign fifo_intf_2278.wr_en = AESL_inst_myproject.layer3_out_925_U.if_write & AESL_inst_myproject.layer3_out_925_U.if_full_n;
    assign fifo_intf_2278.fifo_rd_block = 0;
    assign fifo_intf_2278.fifo_wr_block = 0;
    assign fifo_intf_2278.finish = finish;
    csv_file_dump fifo_csv_dumper_2278;
    csv_file_dump cstatus_csv_dumper_2278;
    df_fifo_monitor fifo_monitor_2278;
    df_fifo_intf fifo_intf_2279(clock,reset);
    assign fifo_intf_2279.rd_en = AESL_inst_myproject.layer3_out_926_U.if_read & AESL_inst_myproject.layer3_out_926_U.if_empty_n;
    assign fifo_intf_2279.wr_en = AESL_inst_myproject.layer3_out_926_U.if_write & AESL_inst_myproject.layer3_out_926_U.if_full_n;
    assign fifo_intf_2279.fifo_rd_block = 0;
    assign fifo_intf_2279.fifo_wr_block = 0;
    assign fifo_intf_2279.finish = finish;
    csv_file_dump fifo_csv_dumper_2279;
    csv_file_dump cstatus_csv_dumper_2279;
    df_fifo_monitor fifo_monitor_2279;
    df_fifo_intf fifo_intf_2280(clock,reset);
    assign fifo_intf_2280.rd_en = AESL_inst_myproject.layer3_out_927_U.if_read & AESL_inst_myproject.layer3_out_927_U.if_empty_n;
    assign fifo_intf_2280.wr_en = AESL_inst_myproject.layer3_out_927_U.if_write & AESL_inst_myproject.layer3_out_927_U.if_full_n;
    assign fifo_intf_2280.fifo_rd_block = 0;
    assign fifo_intf_2280.fifo_wr_block = 0;
    assign fifo_intf_2280.finish = finish;
    csv_file_dump fifo_csv_dumper_2280;
    csv_file_dump cstatus_csv_dumper_2280;
    df_fifo_monitor fifo_monitor_2280;
    df_fifo_intf fifo_intf_2281(clock,reset);
    assign fifo_intf_2281.rd_en = AESL_inst_myproject.layer3_out_928_U.if_read & AESL_inst_myproject.layer3_out_928_U.if_empty_n;
    assign fifo_intf_2281.wr_en = AESL_inst_myproject.layer3_out_928_U.if_write & AESL_inst_myproject.layer3_out_928_U.if_full_n;
    assign fifo_intf_2281.fifo_rd_block = 0;
    assign fifo_intf_2281.fifo_wr_block = 0;
    assign fifo_intf_2281.finish = finish;
    csv_file_dump fifo_csv_dumper_2281;
    csv_file_dump cstatus_csv_dumper_2281;
    df_fifo_monitor fifo_monitor_2281;
    df_fifo_intf fifo_intf_2282(clock,reset);
    assign fifo_intf_2282.rd_en = AESL_inst_myproject.layer3_out_929_U.if_read & AESL_inst_myproject.layer3_out_929_U.if_empty_n;
    assign fifo_intf_2282.wr_en = AESL_inst_myproject.layer3_out_929_U.if_write & AESL_inst_myproject.layer3_out_929_U.if_full_n;
    assign fifo_intf_2282.fifo_rd_block = 0;
    assign fifo_intf_2282.fifo_wr_block = 0;
    assign fifo_intf_2282.finish = finish;
    csv_file_dump fifo_csv_dumper_2282;
    csv_file_dump cstatus_csv_dumper_2282;
    df_fifo_monitor fifo_monitor_2282;
    df_fifo_intf fifo_intf_2283(clock,reset);
    assign fifo_intf_2283.rd_en = AESL_inst_myproject.layer3_out_930_U.if_read & AESL_inst_myproject.layer3_out_930_U.if_empty_n;
    assign fifo_intf_2283.wr_en = AESL_inst_myproject.layer3_out_930_U.if_write & AESL_inst_myproject.layer3_out_930_U.if_full_n;
    assign fifo_intf_2283.fifo_rd_block = 0;
    assign fifo_intf_2283.fifo_wr_block = 0;
    assign fifo_intf_2283.finish = finish;
    csv_file_dump fifo_csv_dumper_2283;
    csv_file_dump cstatus_csv_dumper_2283;
    df_fifo_monitor fifo_monitor_2283;
    df_fifo_intf fifo_intf_2284(clock,reset);
    assign fifo_intf_2284.rd_en = AESL_inst_myproject.layer3_out_931_U.if_read & AESL_inst_myproject.layer3_out_931_U.if_empty_n;
    assign fifo_intf_2284.wr_en = AESL_inst_myproject.layer3_out_931_U.if_write & AESL_inst_myproject.layer3_out_931_U.if_full_n;
    assign fifo_intf_2284.fifo_rd_block = 0;
    assign fifo_intf_2284.fifo_wr_block = 0;
    assign fifo_intf_2284.finish = finish;
    csv_file_dump fifo_csv_dumper_2284;
    csv_file_dump cstatus_csv_dumper_2284;
    df_fifo_monitor fifo_monitor_2284;
    df_fifo_intf fifo_intf_2285(clock,reset);
    assign fifo_intf_2285.rd_en = AESL_inst_myproject.layer3_out_932_U.if_read & AESL_inst_myproject.layer3_out_932_U.if_empty_n;
    assign fifo_intf_2285.wr_en = AESL_inst_myproject.layer3_out_932_U.if_write & AESL_inst_myproject.layer3_out_932_U.if_full_n;
    assign fifo_intf_2285.fifo_rd_block = 0;
    assign fifo_intf_2285.fifo_wr_block = 0;
    assign fifo_intf_2285.finish = finish;
    csv_file_dump fifo_csv_dumper_2285;
    csv_file_dump cstatus_csv_dumper_2285;
    df_fifo_monitor fifo_monitor_2285;
    df_fifo_intf fifo_intf_2286(clock,reset);
    assign fifo_intf_2286.rd_en = AESL_inst_myproject.layer3_out_933_U.if_read & AESL_inst_myproject.layer3_out_933_U.if_empty_n;
    assign fifo_intf_2286.wr_en = AESL_inst_myproject.layer3_out_933_U.if_write & AESL_inst_myproject.layer3_out_933_U.if_full_n;
    assign fifo_intf_2286.fifo_rd_block = 0;
    assign fifo_intf_2286.fifo_wr_block = 0;
    assign fifo_intf_2286.finish = finish;
    csv_file_dump fifo_csv_dumper_2286;
    csv_file_dump cstatus_csv_dumper_2286;
    df_fifo_monitor fifo_monitor_2286;
    df_fifo_intf fifo_intf_2287(clock,reset);
    assign fifo_intf_2287.rd_en = AESL_inst_myproject.layer3_out_934_U.if_read & AESL_inst_myproject.layer3_out_934_U.if_empty_n;
    assign fifo_intf_2287.wr_en = AESL_inst_myproject.layer3_out_934_U.if_write & AESL_inst_myproject.layer3_out_934_U.if_full_n;
    assign fifo_intf_2287.fifo_rd_block = 0;
    assign fifo_intf_2287.fifo_wr_block = 0;
    assign fifo_intf_2287.finish = finish;
    csv_file_dump fifo_csv_dumper_2287;
    csv_file_dump cstatus_csv_dumper_2287;
    df_fifo_monitor fifo_monitor_2287;
    df_fifo_intf fifo_intf_2288(clock,reset);
    assign fifo_intf_2288.rd_en = AESL_inst_myproject.layer3_out_935_U.if_read & AESL_inst_myproject.layer3_out_935_U.if_empty_n;
    assign fifo_intf_2288.wr_en = AESL_inst_myproject.layer3_out_935_U.if_write & AESL_inst_myproject.layer3_out_935_U.if_full_n;
    assign fifo_intf_2288.fifo_rd_block = 0;
    assign fifo_intf_2288.fifo_wr_block = 0;
    assign fifo_intf_2288.finish = finish;
    csv_file_dump fifo_csv_dumper_2288;
    csv_file_dump cstatus_csv_dumper_2288;
    df_fifo_monitor fifo_monitor_2288;
    df_fifo_intf fifo_intf_2289(clock,reset);
    assign fifo_intf_2289.rd_en = AESL_inst_myproject.layer3_out_936_U.if_read & AESL_inst_myproject.layer3_out_936_U.if_empty_n;
    assign fifo_intf_2289.wr_en = AESL_inst_myproject.layer3_out_936_U.if_write & AESL_inst_myproject.layer3_out_936_U.if_full_n;
    assign fifo_intf_2289.fifo_rd_block = 0;
    assign fifo_intf_2289.fifo_wr_block = 0;
    assign fifo_intf_2289.finish = finish;
    csv_file_dump fifo_csv_dumper_2289;
    csv_file_dump cstatus_csv_dumper_2289;
    df_fifo_monitor fifo_monitor_2289;
    df_fifo_intf fifo_intf_2290(clock,reset);
    assign fifo_intf_2290.rd_en = AESL_inst_myproject.layer3_out_937_U.if_read & AESL_inst_myproject.layer3_out_937_U.if_empty_n;
    assign fifo_intf_2290.wr_en = AESL_inst_myproject.layer3_out_937_U.if_write & AESL_inst_myproject.layer3_out_937_U.if_full_n;
    assign fifo_intf_2290.fifo_rd_block = 0;
    assign fifo_intf_2290.fifo_wr_block = 0;
    assign fifo_intf_2290.finish = finish;
    csv_file_dump fifo_csv_dumper_2290;
    csv_file_dump cstatus_csv_dumper_2290;
    df_fifo_monitor fifo_monitor_2290;
    df_fifo_intf fifo_intf_2291(clock,reset);
    assign fifo_intf_2291.rd_en = AESL_inst_myproject.layer3_out_938_U.if_read & AESL_inst_myproject.layer3_out_938_U.if_empty_n;
    assign fifo_intf_2291.wr_en = AESL_inst_myproject.layer3_out_938_U.if_write & AESL_inst_myproject.layer3_out_938_U.if_full_n;
    assign fifo_intf_2291.fifo_rd_block = 0;
    assign fifo_intf_2291.fifo_wr_block = 0;
    assign fifo_intf_2291.finish = finish;
    csv_file_dump fifo_csv_dumper_2291;
    csv_file_dump cstatus_csv_dumper_2291;
    df_fifo_monitor fifo_monitor_2291;
    df_fifo_intf fifo_intf_2292(clock,reset);
    assign fifo_intf_2292.rd_en = AESL_inst_myproject.layer3_out_939_U.if_read & AESL_inst_myproject.layer3_out_939_U.if_empty_n;
    assign fifo_intf_2292.wr_en = AESL_inst_myproject.layer3_out_939_U.if_write & AESL_inst_myproject.layer3_out_939_U.if_full_n;
    assign fifo_intf_2292.fifo_rd_block = 0;
    assign fifo_intf_2292.fifo_wr_block = 0;
    assign fifo_intf_2292.finish = finish;
    csv_file_dump fifo_csv_dumper_2292;
    csv_file_dump cstatus_csv_dumper_2292;
    df_fifo_monitor fifo_monitor_2292;
    df_fifo_intf fifo_intf_2293(clock,reset);
    assign fifo_intf_2293.rd_en = AESL_inst_myproject.layer3_out_940_U.if_read & AESL_inst_myproject.layer3_out_940_U.if_empty_n;
    assign fifo_intf_2293.wr_en = AESL_inst_myproject.layer3_out_940_U.if_write & AESL_inst_myproject.layer3_out_940_U.if_full_n;
    assign fifo_intf_2293.fifo_rd_block = 0;
    assign fifo_intf_2293.fifo_wr_block = 0;
    assign fifo_intf_2293.finish = finish;
    csv_file_dump fifo_csv_dumper_2293;
    csv_file_dump cstatus_csv_dumper_2293;
    df_fifo_monitor fifo_monitor_2293;
    df_fifo_intf fifo_intf_2294(clock,reset);
    assign fifo_intf_2294.rd_en = AESL_inst_myproject.layer3_out_941_U.if_read & AESL_inst_myproject.layer3_out_941_U.if_empty_n;
    assign fifo_intf_2294.wr_en = AESL_inst_myproject.layer3_out_941_U.if_write & AESL_inst_myproject.layer3_out_941_U.if_full_n;
    assign fifo_intf_2294.fifo_rd_block = 0;
    assign fifo_intf_2294.fifo_wr_block = 0;
    assign fifo_intf_2294.finish = finish;
    csv_file_dump fifo_csv_dumper_2294;
    csv_file_dump cstatus_csv_dumper_2294;
    df_fifo_monitor fifo_monitor_2294;
    df_fifo_intf fifo_intf_2295(clock,reset);
    assign fifo_intf_2295.rd_en = AESL_inst_myproject.layer3_out_942_U.if_read & AESL_inst_myproject.layer3_out_942_U.if_empty_n;
    assign fifo_intf_2295.wr_en = AESL_inst_myproject.layer3_out_942_U.if_write & AESL_inst_myproject.layer3_out_942_U.if_full_n;
    assign fifo_intf_2295.fifo_rd_block = 0;
    assign fifo_intf_2295.fifo_wr_block = 0;
    assign fifo_intf_2295.finish = finish;
    csv_file_dump fifo_csv_dumper_2295;
    csv_file_dump cstatus_csv_dumper_2295;
    df_fifo_monitor fifo_monitor_2295;
    df_fifo_intf fifo_intf_2296(clock,reset);
    assign fifo_intf_2296.rd_en = AESL_inst_myproject.layer3_out_943_U.if_read & AESL_inst_myproject.layer3_out_943_U.if_empty_n;
    assign fifo_intf_2296.wr_en = AESL_inst_myproject.layer3_out_943_U.if_write & AESL_inst_myproject.layer3_out_943_U.if_full_n;
    assign fifo_intf_2296.fifo_rd_block = 0;
    assign fifo_intf_2296.fifo_wr_block = 0;
    assign fifo_intf_2296.finish = finish;
    csv_file_dump fifo_csv_dumper_2296;
    csv_file_dump cstatus_csv_dumper_2296;
    df_fifo_monitor fifo_monitor_2296;
    df_fifo_intf fifo_intf_2297(clock,reset);
    assign fifo_intf_2297.rd_en = AESL_inst_myproject.layer3_out_944_U.if_read & AESL_inst_myproject.layer3_out_944_U.if_empty_n;
    assign fifo_intf_2297.wr_en = AESL_inst_myproject.layer3_out_944_U.if_write & AESL_inst_myproject.layer3_out_944_U.if_full_n;
    assign fifo_intf_2297.fifo_rd_block = 0;
    assign fifo_intf_2297.fifo_wr_block = 0;
    assign fifo_intf_2297.finish = finish;
    csv_file_dump fifo_csv_dumper_2297;
    csv_file_dump cstatus_csv_dumper_2297;
    df_fifo_monitor fifo_monitor_2297;
    df_fifo_intf fifo_intf_2298(clock,reset);
    assign fifo_intf_2298.rd_en = AESL_inst_myproject.layer3_out_945_U.if_read & AESL_inst_myproject.layer3_out_945_U.if_empty_n;
    assign fifo_intf_2298.wr_en = AESL_inst_myproject.layer3_out_945_U.if_write & AESL_inst_myproject.layer3_out_945_U.if_full_n;
    assign fifo_intf_2298.fifo_rd_block = 0;
    assign fifo_intf_2298.fifo_wr_block = 0;
    assign fifo_intf_2298.finish = finish;
    csv_file_dump fifo_csv_dumper_2298;
    csv_file_dump cstatus_csv_dumper_2298;
    df_fifo_monitor fifo_monitor_2298;
    df_fifo_intf fifo_intf_2299(clock,reset);
    assign fifo_intf_2299.rd_en = AESL_inst_myproject.layer3_out_946_U.if_read & AESL_inst_myproject.layer3_out_946_U.if_empty_n;
    assign fifo_intf_2299.wr_en = AESL_inst_myproject.layer3_out_946_U.if_write & AESL_inst_myproject.layer3_out_946_U.if_full_n;
    assign fifo_intf_2299.fifo_rd_block = 0;
    assign fifo_intf_2299.fifo_wr_block = 0;
    assign fifo_intf_2299.finish = finish;
    csv_file_dump fifo_csv_dumper_2299;
    csv_file_dump cstatus_csv_dumper_2299;
    df_fifo_monitor fifo_monitor_2299;
    df_fifo_intf fifo_intf_2300(clock,reset);
    assign fifo_intf_2300.rd_en = AESL_inst_myproject.layer3_out_947_U.if_read & AESL_inst_myproject.layer3_out_947_U.if_empty_n;
    assign fifo_intf_2300.wr_en = AESL_inst_myproject.layer3_out_947_U.if_write & AESL_inst_myproject.layer3_out_947_U.if_full_n;
    assign fifo_intf_2300.fifo_rd_block = 0;
    assign fifo_intf_2300.fifo_wr_block = 0;
    assign fifo_intf_2300.finish = finish;
    csv_file_dump fifo_csv_dumper_2300;
    csv_file_dump cstatus_csv_dumper_2300;
    df_fifo_monitor fifo_monitor_2300;
    df_fifo_intf fifo_intf_2301(clock,reset);
    assign fifo_intf_2301.rd_en = AESL_inst_myproject.layer3_out_948_U.if_read & AESL_inst_myproject.layer3_out_948_U.if_empty_n;
    assign fifo_intf_2301.wr_en = AESL_inst_myproject.layer3_out_948_U.if_write & AESL_inst_myproject.layer3_out_948_U.if_full_n;
    assign fifo_intf_2301.fifo_rd_block = 0;
    assign fifo_intf_2301.fifo_wr_block = 0;
    assign fifo_intf_2301.finish = finish;
    csv_file_dump fifo_csv_dumper_2301;
    csv_file_dump cstatus_csv_dumper_2301;
    df_fifo_monitor fifo_monitor_2301;
    df_fifo_intf fifo_intf_2302(clock,reset);
    assign fifo_intf_2302.rd_en = AESL_inst_myproject.layer3_out_949_U.if_read & AESL_inst_myproject.layer3_out_949_U.if_empty_n;
    assign fifo_intf_2302.wr_en = AESL_inst_myproject.layer3_out_949_U.if_write & AESL_inst_myproject.layer3_out_949_U.if_full_n;
    assign fifo_intf_2302.fifo_rd_block = 0;
    assign fifo_intf_2302.fifo_wr_block = 0;
    assign fifo_intf_2302.finish = finish;
    csv_file_dump fifo_csv_dumper_2302;
    csv_file_dump cstatus_csv_dumper_2302;
    df_fifo_monitor fifo_monitor_2302;
    df_fifo_intf fifo_intf_2303(clock,reset);
    assign fifo_intf_2303.rd_en = AESL_inst_myproject.layer3_out_950_U.if_read & AESL_inst_myproject.layer3_out_950_U.if_empty_n;
    assign fifo_intf_2303.wr_en = AESL_inst_myproject.layer3_out_950_U.if_write & AESL_inst_myproject.layer3_out_950_U.if_full_n;
    assign fifo_intf_2303.fifo_rd_block = 0;
    assign fifo_intf_2303.fifo_wr_block = 0;
    assign fifo_intf_2303.finish = finish;
    csv_file_dump fifo_csv_dumper_2303;
    csv_file_dump cstatus_csv_dumper_2303;
    df_fifo_monitor fifo_monitor_2303;
    df_fifo_intf fifo_intf_2304(clock,reset);
    assign fifo_intf_2304.rd_en = AESL_inst_myproject.layer3_out_951_U.if_read & AESL_inst_myproject.layer3_out_951_U.if_empty_n;
    assign fifo_intf_2304.wr_en = AESL_inst_myproject.layer3_out_951_U.if_write & AESL_inst_myproject.layer3_out_951_U.if_full_n;
    assign fifo_intf_2304.fifo_rd_block = 0;
    assign fifo_intf_2304.fifo_wr_block = 0;
    assign fifo_intf_2304.finish = finish;
    csv_file_dump fifo_csv_dumper_2304;
    csv_file_dump cstatus_csv_dumper_2304;
    df_fifo_monitor fifo_monitor_2304;
    df_fifo_intf fifo_intf_2305(clock,reset);
    assign fifo_intf_2305.rd_en = AESL_inst_myproject.layer3_out_952_U.if_read & AESL_inst_myproject.layer3_out_952_U.if_empty_n;
    assign fifo_intf_2305.wr_en = AESL_inst_myproject.layer3_out_952_U.if_write & AESL_inst_myproject.layer3_out_952_U.if_full_n;
    assign fifo_intf_2305.fifo_rd_block = 0;
    assign fifo_intf_2305.fifo_wr_block = 0;
    assign fifo_intf_2305.finish = finish;
    csv_file_dump fifo_csv_dumper_2305;
    csv_file_dump cstatus_csv_dumper_2305;
    df_fifo_monitor fifo_monitor_2305;
    df_fifo_intf fifo_intf_2306(clock,reset);
    assign fifo_intf_2306.rd_en = AESL_inst_myproject.layer3_out_953_U.if_read & AESL_inst_myproject.layer3_out_953_U.if_empty_n;
    assign fifo_intf_2306.wr_en = AESL_inst_myproject.layer3_out_953_U.if_write & AESL_inst_myproject.layer3_out_953_U.if_full_n;
    assign fifo_intf_2306.fifo_rd_block = 0;
    assign fifo_intf_2306.fifo_wr_block = 0;
    assign fifo_intf_2306.finish = finish;
    csv_file_dump fifo_csv_dumper_2306;
    csv_file_dump cstatus_csv_dumper_2306;
    df_fifo_monitor fifo_monitor_2306;
    df_fifo_intf fifo_intf_2307(clock,reset);
    assign fifo_intf_2307.rd_en = AESL_inst_myproject.layer3_out_954_U.if_read & AESL_inst_myproject.layer3_out_954_U.if_empty_n;
    assign fifo_intf_2307.wr_en = AESL_inst_myproject.layer3_out_954_U.if_write & AESL_inst_myproject.layer3_out_954_U.if_full_n;
    assign fifo_intf_2307.fifo_rd_block = 0;
    assign fifo_intf_2307.fifo_wr_block = 0;
    assign fifo_intf_2307.finish = finish;
    csv_file_dump fifo_csv_dumper_2307;
    csv_file_dump cstatus_csv_dumper_2307;
    df_fifo_monitor fifo_monitor_2307;
    df_fifo_intf fifo_intf_2308(clock,reset);
    assign fifo_intf_2308.rd_en = AESL_inst_myproject.layer3_out_955_U.if_read & AESL_inst_myproject.layer3_out_955_U.if_empty_n;
    assign fifo_intf_2308.wr_en = AESL_inst_myproject.layer3_out_955_U.if_write & AESL_inst_myproject.layer3_out_955_U.if_full_n;
    assign fifo_intf_2308.fifo_rd_block = 0;
    assign fifo_intf_2308.fifo_wr_block = 0;
    assign fifo_intf_2308.finish = finish;
    csv_file_dump fifo_csv_dumper_2308;
    csv_file_dump cstatus_csv_dumper_2308;
    df_fifo_monitor fifo_monitor_2308;
    df_fifo_intf fifo_intf_2309(clock,reset);
    assign fifo_intf_2309.rd_en = AESL_inst_myproject.layer3_out_956_U.if_read & AESL_inst_myproject.layer3_out_956_U.if_empty_n;
    assign fifo_intf_2309.wr_en = AESL_inst_myproject.layer3_out_956_U.if_write & AESL_inst_myproject.layer3_out_956_U.if_full_n;
    assign fifo_intf_2309.fifo_rd_block = 0;
    assign fifo_intf_2309.fifo_wr_block = 0;
    assign fifo_intf_2309.finish = finish;
    csv_file_dump fifo_csv_dumper_2309;
    csv_file_dump cstatus_csv_dumper_2309;
    df_fifo_monitor fifo_monitor_2309;
    df_fifo_intf fifo_intf_2310(clock,reset);
    assign fifo_intf_2310.rd_en = AESL_inst_myproject.layer3_out_957_U.if_read & AESL_inst_myproject.layer3_out_957_U.if_empty_n;
    assign fifo_intf_2310.wr_en = AESL_inst_myproject.layer3_out_957_U.if_write & AESL_inst_myproject.layer3_out_957_U.if_full_n;
    assign fifo_intf_2310.fifo_rd_block = 0;
    assign fifo_intf_2310.fifo_wr_block = 0;
    assign fifo_intf_2310.finish = finish;
    csv_file_dump fifo_csv_dumper_2310;
    csv_file_dump cstatus_csv_dumper_2310;
    df_fifo_monitor fifo_monitor_2310;
    df_fifo_intf fifo_intf_2311(clock,reset);
    assign fifo_intf_2311.rd_en = AESL_inst_myproject.layer3_out_958_U.if_read & AESL_inst_myproject.layer3_out_958_U.if_empty_n;
    assign fifo_intf_2311.wr_en = AESL_inst_myproject.layer3_out_958_U.if_write & AESL_inst_myproject.layer3_out_958_U.if_full_n;
    assign fifo_intf_2311.fifo_rd_block = 0;
    assign fifo_intf_2311.fifo_wr_block = 0;
    assign fifo_intf_2311.finish = finish;
    csv_file_dump fifo_csv_dumper_2311;
    csv_file_dump cstatus_csv_dumper_2311;
    df_fifo_monitor fifo_monitor_2311;
    df_fifo_intf fifo_intf_2312(clock,reset);
    assign fifo_intf_2312.rd_en = AESL_inst_myproject.layer3_out_959_U.if_read & AESL_inst_myproject.layer3_out_959_U.if_empty_n;
    assign fifo_intf_2312.wr_en = AESL_inst_myproject.layer3_out_959_U.if_write & AESL_inst_myproject.layer3_out_959_U.if_full_n;
    assign fifo_intf_2312.fifo_rd_block = 0;
    assign fifo_intf_2312.fifo_wr_block = 0;
    assign fifo_intf_2312.finish = finish;
    csv_file_dump fifo_csv_dumper_2312;
    csv_file_dump cstatus_csv_dumper_2312;
    df_fifo_monitor fifo_monitor_2312;
    df_fifo_intf fifo_intf_2313(clock,reset);
    assign fifo_intf_2313.rd_en = AESL_inst_myproject.layer3_out_960_U.if_read & AESL_inst_myproject.layer3_out_960_U.if_empty_n;
    assign fifo_intf_2313.wr_en = AESL_inst_myproject.layer3_out_960_U.if_write & AESL_inst_myproject.layer3_out_960_U.if_full_n;
    assign fifo_intf_2313.fifo_rd_block = 0;
    assign fifo_intf_2313.fifo_wr_block = 0;
    assign fifo_intf_2313.finish = finish;
    csv_file_dump fifo_csv_dumper_2313;
    csv_file_dump cstatus_csv_dumper_2313;
    df_fifo_monitor fifo_monitor_2313;
    df_fifo_intf fifo_intf_2314(clock,reset);
    assign fifo_intf_2314.rd_en = AESL_inst_myproject.layer3_out_961_U.if_read & AESL_inst_myproject.layer3_out_961_U.if_empty_n;
    assign fifo_intf_2314.wr_en = AESL_inst_myproject.layer3_out_961_U.if_write & AESL_inst_myproject.layer3_out_961_U.if_full_n;
    assign fifo_intf_2314.fifo_rd_block = 0;
    assign fifo_intf_2314.fifo_wr_block = 0;
    assign fifo_intf_2314.finish = finish;
    csv_file_dump fifo_csv_dumper_2314;
    csv_file_dump cstatus_csv_dumper_2314;
    df_fifo_monitor fifo_monitor_2314;
    df_fifo_intf fifo_intf_2315(clock,reset);
    assign fifo_intf_2315.rd_en = AESL_inst_myproject.layer3_out_962_U.if_read & AESL_inst_myproject.layer3_out_962_U.if_empty_n;
    assign fifo_intf_2315.wr_en = AESL_inst_myproject.layer3_out_962_U.if_write & AESL_inst_myproject.layer3_out_962_U.if_full_n;
    assign fifo_intf_2315.fifo_rd_block = 0;
    assign fifo_intf_2315.fifo_wr_block = 0;
    assign fifo_intf_2315.finish = finish;
    csv_file_dump fifo_csv_dumper_2315;
    csv_file_dump cstatus_csv_dumper_2315;
    df_fifo_monitor fifo_monitor_2315;
    df_fifo_intf fifo_intf_2316(clock,reset);
    assign fifo_intf_2316.rd_en = AESL_inst_myproject.layer3_out_963_U.if_read & AESL_inst_myproject.layer3_out_963_U.if_empty_n;
    assign fifo_intf_2316.wr_en = AESL_inst_myproject.layer3_out_963_U.if_write & AESL_inst_myproject.layer3_out_963_U.if_full_n;
    assign fifo_intf_2316.fifo_rd_block = 0;
    assign fifo_intf_2316.fifo_wr_block = 0;
    assign fifo_intf_2316.finish = finish;
    csv_file_dump fifo_csv_dumper_2316;
    csv_file_dump cstatus_csv_dumper_2316;
    df_fifo_monitor fifo_monitor_2316;
    df_fifo_intf fifo_intf_2317(clock,reset);
    assign fifo_intf_2317.rd_en = AESL_inst_myproject.layer3_out_964_U.if_read & AESL_inst_myproject.layer3_out_964_U.if_empty_n;
    assign fifo_intf_2317.wr_en = AESL_inst_myproject.layer3_out_964_U.if_write & AESL_inst_myproject.layer3_out_964_U.if_full_n;
    assign fifo_intf_2317.fifo_rd_block = 0;
    assign fifo_intf_2317.fifo_wr_block = 0;
    assign fifo_intf_2317.finish = finish;
    csv_file_dump fifo_csv_dumper_2317;
    csv_file_dump cstatus_csv_dumper_2317;
    df_fifo_monitor fifo_monitor_2317;
    df_fifo_intf fifo_intf_2318(clock,reset);
    assign fifo_intf_2318.rd_en = AESL_inst_myproject.layer3_out_965_U.if_read & AESL_inst_myproject.layer3_out_965_U.if_empty_n;
    assign fifo_intf_2318.wr_en = AESL_inst_myproject.layer3_out_965_U.if_write & AESL_inst_myproject.layer3_out_965_U.if_full_n;
    assign fifo_intf_2318.fifo_rd_block = 0;
    assign fifo_intf_2318.fifo_wr_block = 0;
    assign fifo_intf_2318.finish = finish;
    csv_file_dump fifo_csv_dumper_2318;
    csv_file_dump cstatus_csv_dumper_2318;
    df_fifo_monitor fifo_monitor_2318;
    df_fifo_intf fifo_intf_2319(clock,reset);
    assign fifo_intf_2319.rd_en = AESL_inst_myproject.layer3_out_966_U.if_read & AESL_inst_myproject.layer3_out_966_U.if_empty_n;
    assign fifo_intf_2319.wr_en = AESL_inst_myproject.layer3_out_966_U.if_write & AESL_inst_myproject.layer3_out_966_U.if_full_n;
    assign fifo_intf_2319.fifo_rd_block = 0;
    assign fifo_intf_2319.fifo_wr_block = 0;
    assign fifo_intf_2319.finish = finish;
    csv_file_dump fifo_csv_dumper_2319;
    csv_file_dump cstatus_csv_dumper_2319;
    df_fifo_monitor fifo_monitor_2319;
    df_fifo_intf fifo_intf_2320(clock,reset);
    assign fifo_intf_2320.rd_en = AESL_inst_myproject.layer3_out_967_U.if_read & AESL_inst_myproject.layer3_out_967_U.if_empty_n;
    assign fifo_intf_2320.wr_en = AESL_inst_myproject.layer3_out_967_U.if_write & AESL_inst_myproject.layer3_out_967_U.if_full_n;
    assign fifo_intf_2320.fifo_rd_block = 0;
    assign fifo_intf_2320.fifo_wr_block = 0;
    assign fifo_intf_2320.finish = finish;
    csv_file_dump fifo_csv_dumper_2320;
    csv_file_dump cstatus_csv_dumper_2320;
    df_fifo_monitor fifo_monitor_2320;
    df_fifo_intf fifo_intf_2321(clock,reset);
    assign fifo_intf_2321.rd_en = AESL_inst_myproject.layer3_out_968_U.if_read & AESL_inst_myproject.layer3_out_968_U.if_empty_n;
    assign fifo_intf_2321.wr_en = AESL_inst_myproject.layer3_out_968_U.if_write & AESL_inst_myproject.layer3_out_968_U.if_full_n;
    assign fifo_intf_2321.fifo_rd_block = 0;
    assign fifo_intf_2321.fifo_wr_block = 0;
    assign fifo_intf_2321.finish = finish;
    csv_file_dump fifo_csv_dumper_2321;
    csv_file_dump cstatus_csv_dumper_2321;
    df_fifo_monitor fifo_monitor_2321;
    df_fifo_intf fifo_intf_2322(clock,reset);
    assign fifo_intf_2322.rd_en = AESL_inst_myproject.layer3_out_969_U.if_read & AESL_inst_myproject.layer3_out_969_U.if_empty_n;
    assign fifo_intf_2322.wr_en = AESL_inst_myproject.layer3_out_969_U.if_write & AESL_inst_myproject.layer3_out_969_U.if_full_n;
    assign fifo_intf_2322.fifo_rd_block = 0;
    assign fifo_intf_2322.fifo_wr_block = 0;
    assign fifo_intf_2322.finish = finish;
    csv_file_dump fifo_csv_dumper_2322;
    csv_file_dump cstatus_csv_dumper_2322;
    df_fifo_monitor fifo_monitor_2322;
    df_fifo_intf fifo_intf_2323(clock,reset);
    assign fifo_intf_2323.rd_en = AESL_inst_myproject.layer3_out_970_U.if_read & AESL_inst_myproject.layer3_out_970_U.if_empty_n;
    assign fifo_intf_2323.wr_en = AESL_inst_myproject.layer3_out_970_U.if_write & AESL_inst_myproject.layer3_out_970_U.if_full_n;
    assign fifo_intf_2323.fifo_rd_block = 0;
    assign fifo_intf_2323.fifo_wr_block = 0;
    assign fifo_intf_2323.finish = finish;
    csv_file_dump fifo_csv_dumper_2323;
    csv_file_dump cstatus_csv_dumper_2323;
    df_fifo_monitor fifo_monitor_2323;
    df_fifo_intf fifo_intf_2324(clock,reset);
    assign fifo_intf_2324.rd_en = AESL_inst_myproject.layer3_out_971_U.if_read & AESL_inst_myproject.layer3_out_971_U.if_empty_n;
    assign fifo_intf_2324.wr_en = AESL_inst_myproject.layer3_out_971_U.if_write & AESL_inst_myproject.layer3_out_971_U.if_full_n;
    assign fifo_intf_2324.fifo_rd_block = 0;
    assign fifo_intf_2324.fifo_wr_block = 0;
    assign fifo_intf_2324.finish = finish;
    csv_file_dump fifo_csv_dumper_2324;
    csv_file_dump cstatus_csv_dumper_2324;
    df_fifo_monitor fifo_monitor_2324;
    df_fifo_intf fifo_intf_2325(clock,reset);
    assign fifo_intf_2325.rd_en = AESL_inst_myproject.layer3_out_972_U.if_read & AESL_inst_myproject.layer3_out_972_U.if_empty_n;
    assign fifo_intf_2325.wr_en = AESL_inst_myproject.layer3_out_972_U.if_write & AESL_inst_myproject.layer3_out_972_U.if_full_n;
    assign fifo_intf_2325.fifo_rd_block = 0;
    assign fifo_intf_2325.fifo_wr_block = 0;
    assign fifo_intf_2325.finish = finish;
    csv_file_dump fifo_csv_dumper_2325;
    csv_file_dump cstatus_csv_dumper_2325;
    df_fifo_monitor fifo_monitor_2325;
    df_fifo_intf fifo_intf_2326(clock,reset);
    assign fifo_intf_2326.rd_en = AESL_inst_myproject.layer3_out_973_U.if_read & AESL_inst_myproject.layer3_out_973_U.if_empty_n;
    assign fifo_intf_2326.wr_en = AESL_inst_myproject.layer3_out_973_U.if_write & AESL_inst_myproject.layer3_out_973_U.if_full_n;
    assign fifo_intf_2326.fifo_rd_block = 0;
    assign fifo_intf_2326.fifo_wr_block = 0;
    assign fifo_intf_2326.finish = finish;
    csv_file_dump fifo_csv_dumper_2326;
    csv_file_dump cstatus_csv_dumper_2326;
    df_fifo_monitor fifo_monitor_2326;
    df_fifo_intf fifo_intf_2327(clock,reset);
    assign fifo_intf_2327.rd_en = AESL_inst_myproject.layer3_out_974_U.if_read & AESL_inst_myproject.layer3_out_974_U.if_empty_n;
    assign fifo_intf_2327.wr_en = AESL_inst_myproject.layer3_out_974_U.if_write & AESL_inst_myproject.layer3_out_974_U.if_full_n;
    assign fifo_intf_2327.fifo_rd_block = 0;
    assign fifo_intf_2327.fifo_wr_block = 0;
    assign fifo_intf_2327.finish = finish;
    csv_file_dump fifo_csv_dumper_2327;
    csv_file_dump cstatus_csv_dumper_2327;
    df_fifo_monitor fifo_monitor_2327;
    df_fifo_intf fifo_intf_2328(clock,reset);
    assign fifo_intf_2328.rd_en = AESL_inst_myproject.layer3_out_975_U.if_read & AESL_inst_myproject.layer3_out_975_U.if_empty_n;
    assign fifo_intf_2328.wr_en = AESL_inst_myproject.layer3_out_975_U.if_write & AESL_inst_myproject.layer3_out_975_U.if_full_n;
    assign fifo_intf_2328.fifo_rd_block = 0;
    assign fifo_intf_2328.fifo_wr_block = 0;
    assign fifo_intf_2328.finish = finish;
    csv_file_dump fifo_csv_dumper_2328;
    csv_file_dump cstatus_csv_dumper_2328;
    df_fifo_monitor fifo_monitor_2328;
    df_fifo_intf fifo_intf_2329(clock,reset);
    assign fifo_intf_2329.rd_en = AESL_inst_myproject.layer3_out_976_U.if_read & AESL_inst_myproject.layer3_out_976_U.if_empty_n;
    assign fifo_intf_2329.wr_en = AESL_inst_myproject.layer3_out_976_U.if_write & AESL_inst_myproject.layer3_out_976_U.if_full_n;
    assign fifo_intf_2329.fifo_rd_block = 0;
    assign fifo_intf_2329.fifo_wr_block = 0;
    assign fifo_intf_2329.finish = finish;
    csv_file_dump fifo_csv_dumper_2329;
    csv_file_dump cstatus_csv_dumper_2329;
    df_fifo_monitor fifo_monitor_2329;
    df_fifo_intf fifo_intf_2330(clock,reset);
    assign fifo_intf_2330.rd_en = AESL_inst_myproject.layer3_out_977_U.if_read & AESL_inst_myproject.layer3_out_977_U.if_empty_n;
    assign fifo_intf_2330.wr_en = AESL_inst_myproject.layer3_out_977_U.if_write & AESL_inst_myproject.layer3_out_977_U.if_full_n;
    assign fifo_intf_2330.fifo_rd_block = 0;
    assign fifo_intf_2330.fifo_wr_block = 0;
    assign fifo_intf_2330.finish = finish;
    csv_file_dump fifo_csv_dumper_2330;
    csv_file_dump cstatus_csv_dumper_2330;
    df_fifo_monitor fifo_monitor_2330;
    df_fifo_intf fifo_intf_2331(clock,reset);
    assign fifo_intf_2331.rd_en = AESL_inst_myproject.layer3_out_978_U.if_read & AESL_inst_myproject.layer3_out_978_U.if_empty_n;
    assign fifo_intf_2331.wr_en = AESL_inst_myproject.layer3_out_978_U.if_write & AESL_inst_myproject.layer3_out_978_U.if_full_n;
    assign fifo_intf_2331.fifo_rd_block = 0;
    assign fifo_intf_2331.fifo_wr_block = 0;
    assign fifo_intf_2331.finish = finish;
    csv_file_dump fifo_csv_dumper_2331;
    csv_file_dump cstatus_csv_dumper_2331;
    df_fifo_monitor fifo_monitor_2331;
    df_fifo_intf fifo_intf_2332(clock,reset);
    assign fifo_intf_2332.rd_en = AESL_inst_myproject.layer3_out_979_U.if_read & AESL_inst_myproject.layer3_out_979_U.if_empty_n;
    assign fifo_intf_2332.wr_en = AESL_inst_myproject.layer3_out_979_U.if_write & AESL_inst_myproject.layer3_out_979_U.if_full_n;
    assign fifo_intf_2332.fifo_rd_block = 0;
    assign fifo_intf_2332.fifo_wr_block = 0;
    assign fifo_intf_2332.finish = finish;
    csv_file_dump fifo_csv_dumper_2332;
    csv_file_dump cstatus_csv_dumper_2332;
    df_fifo_monitor fifo_monitor_2332;
    df_fifo_intf fifo_intf_2333(clock,reset);
    assign fifo_intf_2333.rd_en = AESL_inst_myproject.layer3_out_980_U.if_read & AESL_inst_myproject.layer3_out_980_U.if_empty_n;
    assign fifo_intf_2333.wr_en = AESL_inst_myproject.layer3_out_980_U.if_write & AESL_inst_myproject.layer3_out_980_U.if_full_n;
    assign fifo_intf_2333.fifo_rd_block = 0;
    assign fifo_intf_2333.fifo_wr_block = 0;
    assign fifo_intf_2333.finish = finish;
    csv_file_dump fifo_csv_dumper_2333;
    csv_file_dump cstatus_csv_dumper_2333;
    df_fifo_monitor fifo_monitor_2333;
    df_fifo_intf fifo_intf_2334(clock,reset);
    assign fifo_intf_2334.rd_en = AESL_inst_myproject.layer3_out_981_U.if_read & AESL_inst_myproject.layer3_out_981_U.if_empty_n;
    assign fifo_intf_2334.wr_en = AESL_inst_myproject.layer3_out_981_U.if_write & AESL_inst_myproject.layer3_out_981_U.if_full_n;
    assign fifo_intf_2334.fifo_rd_block = 0;
    assign fifo_intf_2334.fifo_wr_block = 0;
    assign fifo_intf_2334.finish = finish;
    csv_file_dump fifo_csv_dumper_2334;
    csv_file_dump cstatus_csv_dumper_2334;
    df_fifo_monitor fifo_monitor_2334;
    df_fifo_intf fifo_intf_2335(clock,reset);
    assign fifo_intf_2335.rd_en = AESL_inst_myproject.layer3_out_982_U.if_read & AESL_inst_myproject.layer3_out_982_U.if_empty_n;
    assign fifo_intf_2335.wr_en = AESL_inst_myproject.layer3_out_982_U.if_write & AESL_inst_myproject.layer3_out_982_U.if_full_n;
    assign fifo_intf_2335.fifo_rd_block = 0;
    assign fifo_intf_2335.fifo_wr_block = 0;
    assign fifo_intf_2335.finish = finish;
    csv_file_dump fifo_csv_dumper_2335;
    csv_file_dump cstatus_csv_dumper_2335;
    df_fifo_monitor fifo_monitor_2335;
    df_fifo_intf fifo_intf_2336(clock,reset);
    assign fifo_intf_2336.rd_en = AESL_inst_myproject.layer3_out_983_U.if_read & AESL_inst_myproject.layer3_out_983_U.if_empty_n;
    assign fifo_intf_2336.wr_en = AESL_inst_myproject.layer3_out_983_U.if_write & AESL_inst_myproject.layer3_out_983_U.if_full_n;
    assign fifo_intf_2336.fifo_rd_block = 0;
    assign fifo_intf_2336.fifo_wr_block = 0;
    assign fifo_intf_2336.finish = finish;
    csv_file_dump fifo_csv_dumper_2336;
    csv_file_dump cstatus_csv_dumper_2336;
    df_fifo_monitor fifo_monitor_2336;
    df_fifo_intf fifo_intf_2337(clock,reset);
    assign fifo_intf_2337.rd_en = AESL_inst_myproject.layer3_out_984_U.if_read & AESL_inst_myproject.layer3_out_984_U.if_empty_n;
    assign fifo_intf_2337.wr_en = AESL_inst_myproject.layer3_out_984_U.if_write & AESL_inst_myproject.layer3_out_984_U.if_full_n;
    assign fifo_intf_2337.fifo_rd_block = 0;
    assign fifo_intf_2337.fifo_wr_block = 0;
    assign fifo_intf_2337.finish = finish;
    csv_file_dump fifo_csv_dumper_2337;
    csv_file_dump cstatus_csv_dumper_2337;
    df_fifo_monitor fifo_monitor_2337;
    df_fifo_intf fifo_intf_2338(clock,reset);
    assign fifo_intf_2338.rd_en = AESL_inst_myproject.layer3_out_985_U.if_read & AESL_inst_myproject.layer3_out_985_U.if_empty_n;
    assign fifo_intf_2338.wr_en = AESL_inst_myproject.layer3_out_985_U.if_write & AESL_inst_myproject.layer3_out_985_U.if_full_n;
    assign fifo_intf_2338.fifo_rd_block = 0;
    assign fifo_intf_2338.fifo_wr_block = 0;
    assign fifo_intf_2338.finish = finish;
    csv_file_dump fifo_csv_dumper_2338;
    csv_file_dump cstatus_csv_dumper_2338;
    df_fifo_monitor fifo_monitor_2338;
    df_fifo_intf fifo_intf_2339(clock,reset);
    assign fifo_intf_2339.rd_en = AESL_inst_myproject.layer3_out_986_U.if_read & AESL_inst_myproject.layer3_out_986_U.if_empty_n;
    assign fifo_intf_2339.wr_en = AESL_inst_myproject.layer3_out_986_U.if_write & AESL_inst_myproject.layer3_out_986_U.if_full_n;
    assign fifo_intf_2339.fifo_rd_block = 0;
    assign fifo_intf_2339.fifo_wr_block = 0;
    assign fifo_intf_2339.finish = finish;
    csv_file_dump fifo_csv_dumper_2339;
    csv_file_dump cstatus_csv_dumper_2339;
    df_fifo_monitor fifo_monitor_2339;
    df_fifo_intf fifo_intf_2340(clock,reset);
    assign fifo_intf_2340.rd_en = AESL_inst_myproject.layer3_out_987_U.if_read & AESL_inst_myproject.layer3_out_987_U.if_empty_n;
    assign fifo_intf_2340.wr_en = AESL_inst_myproject.layer3_out_987_U.if_write & AESL_inst_myproject.layer3_out_987_U.if_full_n;
    assign fifo_intf_2340.fifo_rd_block = 0;
    assign fifo_intf_2340.fifo_wr_block = 0;
    assign fifo_intf_2340.finish = finish;
    csv_file_dump fifo_csv_dumper_2340;
    csv_file_dump cstatus_csv_dumper_2340;
    df_fifo_monitor fifo_monitor_2340;
    df_fifo_intf fifo_intf_2341(clock,reset);
    assign fifo_intf_2341.rd_en = AESL_inst_myproject.layer3_out_988_U.if_read & AESL_inst_myproject.layer3_out_988_U.if_empty_n;
    assign fifo_intf_2341.wr_en = AESL_inst_myproject.layer3_out_988_U.if_write & AESL_inst_myproject.layer3_out_988_U.if_full_n;
    assign fifo_intf_2341.fifo_rd_block = 0;
    assign fifo_intf_2341.fifo_wr_block = 0;
    assign fifo_intf_2341.finish = finish;
    csv_file_dump fifo_csv_dumper_2341;
    csv_file_dump cstatus_csv_dumper_2341;
    df_fifo_monitor fifo_monitor_2341;
    df_fifo_intf fifo_intf_2342(clock,reset);
    assign fifo_intf_2342.rd_en = AESL_inst_myproject.layer3_out_989_U.if_read & AESL_inst_myproject.layer3_out_989_U.if_empty_n;
    assign fifo_intf_2342.wr_en = AESL_inst_myproject.layer3_out_989_U.if_write & AESL_inst_myproject.layer3_out_989_U.if_full_n;
    assign fifo_intf_2342.fifo_rd_block = 0;
    assign fifo_intf_2342.fifo_wr_block = 0;
    assign fifo_intf_2342.finish = finish;
    csv_file_dump fifo_csv_dumper_2342;
    csv_file_dump cstatus_csv_dumper_2342;
    df_fifo_monitor fifo_monitor_2342;
    df_fifo_intf fifo_intf_2343(clock,reset);
    assign fifo_intf_2343.rd_en = AESL_inst_myproject.layer3_out_990_U.if_read & AESL_inst_myproject.layer3_out_990_U.if_empty_n;
    assign fifo_intf_2343.wr_en = AESL_inst_myproject.layer3_out_990_U.if_write & AESL_inst_myproject.layer3_out_990_U.if_full_n;
    assign fifo_intf_2343.fifo_rd_block = 0;
    assign fifo_intf_2343.fifo_wr_block = 0;
    assign fifo_intf_2343.finish = finish;
    csv_file_dump fifo_csv_dumper_2343;
    csv_file_dump cstatus_csv_dumper_2343;
    df_fifo_monitor fifo_monitor_2343;
    df_fifo_intf fifo_intf_2344(clock,reset);
    assign fifo_intf_2344.rd_en = AESL_inst_myproject.layer3_out_991_U.if_read & AESL_inst_myproject.layer3_out_991_U.if_empty_n;
    assign fifo_intf_2344.wr_en = AESL_inst_myproject.layer3_out_991_U.if_write & AESL_inst_myproject.layer3_out_991_U.if_full_n;
    assign fifo_intf_2344.fifo_rd_block = 0;
    assign fifo_intf_2344.fifo_wr_block = 0;
    assign fifo_intf_2344.finish = finish;
    csv_file_dump fifo_csv_dumper_2344;
    csv_file_dump cstatus_csv_dumper_2344;
    df_fifo_monitor fifo_monitor_2344;
    df_fifo_intf fifo_intf_2345(clock,reset);
    assign fifo_intf_2345.rd_en = AESL_inst_myproject.layer3_out_992_U.if_read & AESL_inst_myproject.layer3_out_992_U.if_empty_n;
    assign fifo_intf_2345.wr_en = AESL_inst_myproject.layer3_out_992_U.if_write & AESL_inst_myproject.layer3_out_992_U.if_full_n;
    assign fifo_intf_2345.fifo_rd_block = 0;
    assign fifo_intf_2345.fifo_wr_block = 0;
    assign fifo_intf_2345.finish = finish;
    csv_file_dump fifo_csv_dumper_2345;
    csv_file_dump cstatus_csv_dumper_2345;
    df_fifo_monitor fifo_monitor_2345;
    df_fifo_intf fifo_intf_2346(clock,reset);
    assign fifo_intf_2346.rd_en = AESL_inst_myproject.layer3_out_993_U.if_read & AESL_inst_myproject.layer3_out_993_U.if_empty_n;
    assign fifo_intf_2346.wr_en = AESL_inst_myproject.layer3_out_993_U.if_write & AESL_inst_myproject.layer3_out_993_U.if_full_n;
    assign fifo_intf_2346.fifo_rd_block = 0;
    assign fifo_intf_2346.fifo_wr_block = 0;
    assign fifo_intf_2346.finish = finish;
    csv_file_dump fifo_csv_dumper_2346;
    csv_file_dump cstatus_csv_dumper_2346;
    df_fifo_monitor fifo_monitor_2346;
    df_fifo_intf fifo_intf_2347(clock,reset);
    assign fifo_intf_2347.rd_en = AESL_inst_myproject.layer3_out_994_U.if_read & AESL_inst_myproject.layer3_out_994_U.if_empty_n;
    assign fifo_intf_2347.wr_en = AESL_inst_myproject.layer3_out_994_U.if_write & AESL_inst_myproject.layer3_out_994_U.if_full_n;
    assign fifo_intf_2347.fifo_rd_block = 0;
    assign fifo_intf_2347.fifo_wr_block = 0;
    assign fifo_intf_2347.finish = finish;
    csv_file_dump fifo_csv_dumper_2347;
    csv_file_dump cstatus_csv_dumper_2347;
    df_fifo_monitor fifo_monitor_2347;
    df_fifo_intf fifo_intf_2348(clock,reset);
    assign fifo_intf_2348.rd_en = AESL_inst_myproject.layer3_out_995_U.if_read & AESL_inst_myproject.layer3_out_995_U.if_empty_n;
    assign fifo_intf_2348.wr_en = AESL_inst_myproject.layer3_out_995_U.if_write & AESL_inst_myproject.layer3_out_995_U.if_full_n;
    assign fifo_intf_2348.fifo_rd_block = 0;
    assign fifo_intf_2348.fifo_wr_block = 0;
    assign fifo_intf_2348.finish = finish;
    csv_file_dump fifo_csv_dumper_2348;
    csv_file_dump cstatus_csv_dumper_2348;
    df_fifo_monitor fifo_monitor_2348;
    df_fifo_intf fifo_intf_2349(clock,reset);
    assign fifo_intf_2349.rd_en = AESL_inst_myproject.layer3_out_996_U.if_read & AESL_inst_myproject.layer3_out_996_U.if_empty_n;
    assign fifo_intf_2349.wr_en = AESL_inst_myproject.layer3_out_996_U.if_write & AESL_inst_myproject.layer3_out_996_U.if_full_n;
    assign fifo_intf_2349.fifo_rd_block = 0;
    assign fifo_intf_2349.fifo_wr_block = 0;
    assign fifo_intf_2349.finish = finish;
    csv_file_dump fifo_csv_dumper_2349;
    csv_file_dump cstatus_csv_dumper_2349;
    df_fifo_monitor fifo_monitor_2349;
    df_fifo_intf fifo_intf_2350(clock,reset);
    assign fifo_intf_2350.rd_en = AESL_inst_myproject.layer3_out_997_U.if_read & AESL_inst_myproject.layer3_out_997_U.if_empty_n;
    assign fifo_intf_2350.wr_en = AESL_inst_myproject.layer3_out_997_U.if_write & AESL_inst_myproject.layer3_out_997_U.if_full_n;
    assign fifo_intf_2350.fifo_rd_block = 0;
    assign fifo_intf_2350.fifo_wr_block = 0;
    assign fifo_intf_2350.finish = finish;
    csv_file_dump fifo_csv_dumper_2350;
    csv_file_dump cstatus_csv_dumper_2350;
    df_fifo_monitor fifo_monitor_2350;
    df_fifo_intf fifo_intf_2351(clock,reset);
    assign fifo_intf_2351.rd_en = AESL_inst_myproject.layer3_out_998_U.if_read & AESL_inst_myproject.layer3_out_998_U.if_empty_n;
    assign fifo_intf_2351.wr_en = AESL_inst_myproject.layer3_out_998_U.if_write & AESL_inst_myproject.layer3_out_998_U.if_full_n;
    assign fifo_intf_2351.fifo_rd_block = 0;
    assign fifo_intf_2351.fifo_wr_block = 0;
    assign fifo_intf_2351.finish = finish;
    csv_file_dump fifo_csv_dumper_2351;
    csv_file_dump cstatus_csv_dumper_2351;
    df_fifo_monitor fifo_monitor_2351;
    df_fifo_intf fifo_intf_2352(clock,reset);
    assign fifo_intf_2352.rd_en = AESL_inst_myproject.layer3_out_999_U.if_read & AESL_inst_myproject.layer3_out_999_U.if_empty_n;
    assign fifo_intf_2352.wr_en = AESL_inst_myproject.layer3_out_999_U.if_write & AESL_inst_myproject.layer3_out_999_U.if_full_n;
    assign fifo_intf_2352.fifo_rd_block = 0;
    assign fifo_intf_2352.fifo_wr_block = 0;
    assign fifo_intf_2352.finish = finish;
    csv_file_dump fifo_csv_dumper_2352;
    csv_file_dump cstatus_csv_dumper_2352;
    df_fifo_monitor fifo_monitor_2352;
    df_fifo_intf fifo_intf_2353(clock,reset);
    assign fifo_intf_2353.rd_en = AESL_inst_myproject.layer3_out_1000_U.if_read & AESL_inst_myproject.layer3_out_1000_U.if_empty_n;
    assign fifo_intf_2353.wr_en = AESL_inst_myproject.layer3_out_1000_U.if_write & AESL_inst_myproject.layer3_out_1000_U.if_full_n;
    assign fifo_intf_2353.fifo_rd_block = 0;
    assign fifo_intf_2353.fifo_wr_block = 0;
    assign fifo_intf_2353.finish = finish;
    csv_file_dump fifo_csv_dumper_2353;
    csv_file_dump cstatus_csv_dumper_2353;
    df_fifo_monitor fifo_monitor_2353;
    df_fifo_intf fifo_intf_2354(clock,reset);
    assign fifo_intf_2354.rd_en = AESL_inst_myproject.layer3_out_1001_U.if_read & AESL_inst_myproject.layer3_out_1001_U.if_empty_n;
    assign fifo_intf_2354.wr_en = AESL_inst_myproject.layer3_out_1001_U.if_write & AESL_inst_myproject.layer3_out_1001_U.if_full_n;
    assign fifo_intf_2354.fifo_rd_block = 0;
    assign fifo_intf_2354.fifo_wr_block = 0;
    assign fifo_intf_2354.finish = finish;
    csv_file_dump fifo_csv_dumper_2354;
    csv_file_dump cstatus_csv_dumper_2354;
    df_fifo_monitor fifo_monitor_2354;
    df_fifo_intf fifo_intf_2355(clock,reset);
    assign fifo_intf_2355.rd_en = AESL_inst_myproject.layer3_out_1002_U.if_read & AESL_inst_myproject.layer3_out_1002_U.if_empty_n;
    assign fifo_intf_2355.wr_en = AESL_inst_myproject.layer3_out_1002_U.if_write & AESL_inst_myproject.layer3_out_1002_U.if_full_n;
    assign fifo_intf_2355.fifo_rd_block = 0;
    assign fifo_intf_2355.fifo_wr_block = 0;
    assign fifo_intf_2355.finish = finish;
    csv_file_dump fifo_csv_dumper_2355;
    csv_file_dump cstatus_csv_dumper_2355;
    df_fifo_monitor fifo_monitor_2355;
    df_fifo_intf fifo_intf_2356(clock,reset);
    assign fifo_intf_2356.rd_en = AESL_inst_myproject.layer3_out_1003_U.if_read & AESL_inst_myproject.layer3_out_1003_U.if_empty_n;
    assign fifo_intf_2356.wr_en = AESL_inst_myproject.layer3_out_1003_U.if_write & AESL_inst_myproject.layer3_out_1003_U.if_full_n;
    assign fifo_intf_2356.fifo_rd_block = 0;
    assign fifo_intf_2356.fifo_wr_block = 0;
    assign fifo_intf_2356.finish = finish;
    csv_file_dump fifo_csv_dumper_2356;
    csv_file_dump cstatus_csv_dumper_2356;
    df_fifo_monitor fifo_monitor_2356;
    df_fifo_intf fifo_intf_2357(clock,reset);
    assign fifo_intf_2357.rd_en = AESL_inst_myproject.layer3_out_1004_U.if_read & AESL_inst_myproject.layer3_out_1004_U.if_empty_n;
    assign fifo_intf_2357.wr_en = AESL_inst_myproject.layer3_out_1004_U.if_write & AESL_inst_myproject.layer3_out_1004_U.if_full_n;
    assign fifo_intf_2357.fifo_rd_block = 0;
    assign fifo_intf_2357.fifo_wr_block = 0;
    assign fifo_intf_2357.finish = finish;
    csv_file_dump fifo_csv_dumper_2357;
    csv_file_dump cstatus_csv_dumper_2357;
    df_fifo_monitor fifo_monitor_2357;
    df_fifo_intf fifo_intf_2358(clock,reset);
    assign fifo_intf_2358.rd_en = AESL_inst_myproject.layer3_out_1005_U.if_read & AESL_inst_myproject.layer3_out_1005_U.if_empty_n;
    assign fifo_intf_2358.wr_en = AESL_inst_myproject.layer3_out_1005_U.if_write & AESL_inst_myproject.layer3_out_1005_U.if_full_n;
    assign fifo_intf_2358.fifo_rd_block = 0;
    assign fifo_intf_2358.fifo_wr_block = 0;
    assign fifo_intf_2358.finish = finish;
    csv_file_dump fifo_csv_dumper_2358;
    csv_file_dump cstatus_csv_dumper_2358;
    df_fifo_monitor fifo_monitor_2358;
    df_fifo_intf fifo_intf_2359(clock,reset);
    assign fifo_intf_2359.rd_en = AESL_inst_myproject.layer3_out_1006_U.if_read & AESL_inst_myproject.layer3_out_1006_U.if_empty_n;
    assign fifo_intf_2359.wr_en = AESL_inst_myproject.layer3_out_1006_U.if_write & AESL_inst_myproject.layer3_out_1006_U.if_full_n;
    assign fifo_intf_2359.fifo_rd_block = 0;
    assign fifo_intf_2359.fifo_wr_block = 0;
    assign fifo_intf_2359.finish = finish;
    csv_file_dump fifo_csv_dumper_2359;
    csv_file_dump cstatus_csv_dumper_2359;
    df_fifo_monitor fifo_monitor_2359;
    df_fifo_intf fifo_intf_2360(clock,reset);
    assign fifo_intf_2360.rd_en = AESL_inst_myproject.layer3_out_1007_U.if_read & AESL_inst_myproject.layer3_out_1007_U.if_empty_n;
    assign fifo_intf_2360.wr_en = AESL_inst_myproject.layer3_out_1007_U.if_write & AESL_inst_myproject.layer3_out_1007_U.if_full_n;
    assign fifo_intf_2360.fifo_rd_block = 0;
    assign fifo_intf_2360.fifo_wr_block = 0;
    assign fifo_intf_2360.finish = finish;
    csv_file_dump fifo_csv_dumper_2360;
    csv_file_dump cstatus_csv_dumper_2360;
    df_fifo_monitor fifo_monitor_2360;
    df_fifo_intf fifo_intf_2361(clock,reset);
    assign fifo_intf_2361.rd_en = AESL_inst_myproject.layer3_out_1008_U.if_read & AESL_inst_myproject.layer3_out_1008_U.if_empty_n;
    assign fifo_intf_2361.wr_en = AESL_inst_myproject.layer3_out_1008_U.if_write & AESL_inst_myproject.layer3_out_1008_U.if_full_n;
    assign fifo_intf_2361.fifo_rd_block = 0;
    assign fifo_intf_2361.fifo_wr_block = 0;
    assign fifo_intf_2361.finish = finish;
    csv_file_dump fifo_csv_dumper_2361;
    csv_file_dump cstatus_csv_dumper_2361;
    df_fifo_monitor fifo_monitor_2361;
    df_fifo_intf fifo_intf_2362(clock,reset);
    assign fifo_intf_2362.rd_en = AESL_inst_myproject.layer3_out_1009_U.if_read & AESL_inst_myproject.layer3_out_1009_U.if_empty_n;
    assign fifo_intf_2362.wr_en = AESL_inst_myproject.layer3_out_1009_U.if_write & AESL_inst_myproject.layer3_out_1009_U.if_full_n;
    assign fifo_intf_2362.fifo_rd_block = 0;
    assign fifo_intf_2362.fifo_wr_block = 0;
    assign fifo_intf_2362.finish = finish;
    csv_file_dump fifo_csv_dumper_2362;
    csv_file_dump cstatus_csv_dumper_2362;
    df_fifo_monitor fifo_monitor_2362;
    df_fifo_intf fifo_intf_2363(clock,reset);
    assign fifo_intf_2363.rd_en = AESL_inst_myproject.layer3_out_1010_U.if_read & AESL_inst_myproject.layer3_out_1010_U.if_empty_n;
    assign fifo_intf_2363.wr_en = AESL_inst_myproject.layer3_out_1010_U.if_write & AESL_inst_myproject.layer3_out_1010_U.if_full_n;
    assign fifo_intf_2363.fifo_rd_block = 0;
    assign fifo_intf_2363.fifo_wr_block = 0;
    assign fifo_intf_2363.finish = finish;
    csv_file_dump fifo_csv_dumper_2363;
    csv_file_dump cstatus_csv_dumper_2363;
    df_fifo_monitor fifo_monitor_2363;
    df_fifo_intf fifo_intf_2364(clock,reset);
    assign fifo_intf_2364.rd_en = AESL_inst_myproject.layer3_out_1011_U.if_read & AESL_inst_myproject.layer3_out_1011_U.if_empty_n;
    assign fifo_intf_2364.wr_en = AESL_inst_myproject.layer3_out_1011_U.if_write & AESL_inst_myproject.layer3_out_1011_U.if_full_n;
    assign fifo_intf_2364.fifo_rd_block = 0;
    assign fifo_intf_2364.fifo_wr_block = 0;
    assign fifo_intf_2364.finish = finish;
    csv_file_dump fifo_csv_dumper_2364;
    csv_file_dump cstatus_csv_dumper_2364;
    df_fifo_monitor fifo_monitor_2364;
    df_fifo_intf fifo_intf_2365(clock,reset);
    assign fifo_intf_2365.rd_en = AESL_inst_myproject.layer3_out_1012_U.if_read & AESL_inst_myproject.layer3_out_1012_U.if_empty_n;
    assign fifo_intf_2365.wr_en = AESL_inst_myproject.layer3_out_1012_U.if_write & AESL_inst_myproject.layer3_out_1012_U.if_full_n;
    assign fifo_intf_2365.fifo_rd_block = 0;
    assign fifo_intf_2365.fifo_wr_block = 0;
    assign fifo_intf_2365.finish = finish;
    csv_file_dump fifo_csv_dumper_2365;
    csv_file_dump cstatus_csv_dumper_2365;
    df_fifo_monitor fifo_monitor_2365;
    df_fifo_intf fifo_intf_2366(clock,reset);
    assign fifo_intf_2366.rd_en = AESL_inst_myproject.layer3_out_1013_U.if_read & AESL_inst_myproject.layer3_out_1013_U.if_empty_n;
    assign fifo_intf_2366.wr_en = AESL_inst_myproject.layer3_out_1013_U.if_write & AESL_inst_myproject.layer3_out_1013_U.if_full_n;
    assign fifo_intf_2366.fifo_rd_block = 0;
    assign fifo_intf_2366.fifo_wr_block = 0;
    assign fifo_intf_2366.finish = finish;
    csv_file_dump fifo_csv_dumper_2366;
    csv_file_dump cstatus_csv_dumper_2366;
    df_fifo_monitor fifo_monitor_2366;
    df_fifo_intf fifo_intf_2367(clock,reset);
    assign fifo_intf_2367.rd_en = AESL_inst_myproject.layer3_out_1014_U.if_read & AESL_inst_myproject.layer3_out_1014_U.if_empty_n;
    assign fifo_intf_2367.wr_en = AESL_inst_myproject.layer3_out_1014_U.if_write & AESL_inst_myproject.layer3_out_1014_U.if_full_n;
    assign fifo_intf_2367.fifo_rd_block = 0;
    assign fifo_intf_2367.fifo_wr_block = 0;
    assign fifo_intf_2367.finish = finish;
    csv_file_dump fifo_csv_dumper_2367;
    csv_file_dump cstatus_csv_dumper_2367;
    df_fifo_monitor fifo_monitor_2367;
    df_fifo_intf fifo_intf_2368(clock,reset);
    assign fifo_intf_2368.rd_en = AESL_inst_myproject.layer3_out_1015_U.if_read & AESL_inst_myproject.layer3_out_1015_U.if_empty_n;
    assign fifo_intf_2368.wr_en = AESL_inst_myproject.layer3_out_1015_U.if_write & AESL_inst_myproject.layer3_out_1015_U.if_full_n;
    assign fifo_intf_2368.fifo_rd_block = 0;
    assign fifo_intf_2368.fifo_wr_block = 0;
    assign fifo_intf_2368.finish = finish;
    csv_file_dump fifo_csv_dumper_2368;
    csv_file_dump cstatus_csv_dumper_2368;
    df_fifo_monitor fifo_monitor_2368;
    df_fifo_intf fifo_intf_2369(clock,reset);
    assign fifo_intf_2369.rd_en = AESL_inst_myproject.layer3_out_1016_U.if_read & AESL_inst_myproject.layer3_out_1016_U.if_empty_n;
    assign fifo_intf_2369.wr_en = AESL_inst_myproject.layer3_out_1016_U.if_write & AESL_inst_myproject.layer3_out_1016_U.if_full_n;
    assign fifo_intf_2369.fifo_rd_block = 0;
    assign fifo_intf_2369.fifo_wr_block = 0;
    assign fifo_intf_2369.finish = finish;
    csv_file_dump fifo_csv_dumper_2369;
    csv_file_dump cstatus_csv_dumper_2369;
    df_fifo_monitor fifo_monitor_2369;
    df_fifo_intf fifo_intf_2370(clock,reset);
    assign fifo_intf_2370.rd_en = AESL_inst_myproject.layer3_out_1017_U.if_read & AESL_inst_myproject.layer3_out_1017_U.if_empty_n;
    assign fifo_intf_2370.wr_en = AESL_inst_myproject.layer3_out_1017_U.if_write & AESL_inst_myproject.layer3_out_1017_U.if_full_n;
    assign fifo_intf_2370.fifo_rd_block = 0;
    assign fifo_intf_2370.fifo_wr_block = 0;
    assign fifo_intf_2370.finish = finish;
    csv_file_dump fifo_csv_dumper_2370;
    csv_file_dump cstatus_csv_dumper_2370;
    df_fifo_monitor fifo_monitor_2370;
    df_fifo_intf fifo_intf_2371(clock,reset);
    assign fifo_intf_2371.rd_en = AESL_inst_myproject.layer3_out_1018_U.if_read & AESL_inst_myproject.layer3_out_1018_U.if_empty_n;
    assign fifo_intf_2371.wr_en = AESL_inst_myproject.layer3_out_1018_U.if_write & AESL_inst_myproject.layer3_out_1018_U.if_full_n;
    assign fifo_intf_2371.fifo_rd_block = 0;
    assign fifo_intf_2371.fifo_wr_block = 0;
    assign fifo_intf_2371.finish = finish;
    csv_file_dump fifo_csv_dumper_2371;
    csv_file_dump cstatus_csv_dumper_2371;
    df_fifo_monitor fifo_monitor_2371;
    df_fifo_intf fifo_intf_2372(clock,reset);
    assign fifo_intf_2372.rd_en = AESL_inst_myproject.layer3_out_1019_U.if_read & AESL_inst_myproject.layer3_out_1019_U.if_empty_n;
    assign fifo_intf_2372.wr_en = AESL_inst_myproject.layer3_out_1019_U.if_write & AESL_inst_myproject.layer3_out_1019_U.if_full_n;
    assign fifo_intf_2372.fifo_rd_block = 0;
    assign fifo_intf_2372.fifo_wr_block = 0;
    assign fifo_intf_2372.finish = finish;
    csv_file_dump fifo_csv_dumper_2372;
    csv_file_dump cstatus_csv_dumper_2372;
    df_fifo_monitor fifo_monitor_2372;
    df_fifo_intf fifo_intf_2373(clock,reset);
    assign fifo_intf_2373.rd_en = AESL_inst_myproject.layer3_out_1020_U.if_read & AESL_inst_myproject.layer3_out_1020_U.if_empty_n;
    assign fifo_intf_2373.wr_en = AESL_inst_myproject.layer3_out_1020_U.if_write & AESL_inst_myproject.layer3_out_1020_U.if_full_n;
    assign fifo_intf_2373.fifo_rd_block = 0;
    assign fifo_intf_2373.fifo_wr_block = 0;
    assign fifo_intf_2373.finish = finish;
    csv_file_dump fifo_csv_dumper_2373;
    csv_file_dump cstatus_csv_dumper_2373;
    df_fifo_monitor fifo_monitor_2373;
    df_fifo_intf fifo_intf_2374(clock,reset);
    assign fifo_intf_2374.rd_en = AESL_inst_myproject.layer3_out_1021_U.if_read & AESL_inst_myproject.layer3_out_1021_U.if_empty_n;
    assign fifo_intf_2374.wr_en = AESL_inst_myproject.layer3_out_1021_U.if_write & AESL_inst_myproject.layer3_out_1021_U.if_full_n;
    assign fifo_intf_2374.fifo_rd_block = 0;
    assign fifo_intf_2374.fifo_wr_block = 0;
    assign fifo_intf_2374.finish = finish;
    csv_file_dump fifo_csv_dumper_2374;
    csv_file_dump cstatus_csv_dumper_2374;
    df_fifo_monitor fifo_monitor_2374;
    df_fifo_intf fifo_intf_2375(clock,reset);
    assign fifo_intf_2375.rd_en = AESL_inst_myproject.layer3_out_1022_U.if_read & AESL_inst_myproject.layer3_out_1022_U.if_empty_n;
    assign fifo_intf_2375.wr_en = AESL_inst_myproject.layer3_out_1022_U.if_write & AESL_inst_myproject.layer3_out_1022_U.if_full_n;
    assign fifo_intf_2375.fifo_rd_block = 0;
    assign fifo_intf_2375.fifo_wr_block = 0;
    assign fifo_intf_2375.finish = finish;
    csv_file_dump fifo_csv_dumper_2375;
    csv_file_dump cstatus_csv_dumper_2375;
    df_fifo_monitor fifo_monitor_2375;
    df_fifo_intf fifo_intf_2376(clock,reset);
    assign fifo_intf_2376.rd_en = AESL_inst_myproject.layer3_out_1023_U.if_read & AESL_inst_myproject.layer3_out_1023_U.if_empty_n;
    assign fifo_intf_2376.wr_en = AESL_inst_myproject.layer3_out_1023_U.if_write & AESL_inst_myproject.layer3_out_1023_U.if_full_n;
    assign fifo_intf_2376.fifo_rd_block = 0;
    assign fifo_intf_2376.fifo_wr_block = 0;
    assign fifo_intf_2376.finish = finish;
    csv_file_dump fifo_csv_dumper_2376;
    csv_file_dump cstatus_csv_dumper_2376;
    df_fifo_monitor fifo_monitor_2376;
    df_fifo_intf fifo_intf_2377(clock,reset);
    assign fifo_intf_2377.rd_en = AESL_inst_myproject.layer3_out_1024_U.if_read & AESL_inst_myproject.layer3_out_1024_U.if_empty_n;
    assign fifo_intf_2377.wr_en = AESL_inst_myproject.layer3_out_1024_U.if_write & AESL_inst_myproject.layer3_out_1024_U.if_full_n;
    assign fifo_intf_2377.fifo_rd_block = 0;
    assign fifo_intf_2377.fifo_wr_block = 0;
    assign fifo_intf_2377.finish = finish;
    csv_file_dump fifo_csv_dumper_2377;
    csv_file_dump cstatus_csv_dumper_2377;
    df_fifo_monitor fifo_monitor_2377;
    df_fifo_intf fifo_intf_2378(clock,reset);
    assign fifo_intf_2378.rd_en = AESL_inst_myproject.layer3_out_1025_U.if_read & AESL_inst_myproject.layer3_out_1025_U.if_empty_n;
    assign fifo_intf_2378.wr_en = AESL_inst_myproject.layer3_out_1025_U.if_write & AESL_inst_myproject.layer3_out_1025_U.if_full_n;
    assign fifo_intf_2378.fifo_rd_block = 0;
    assign fifo_intf_2378.fifo_wr_block = 0;
    assign fifo_intf_2378.finish = finish;
    csv_file_dump fifo_csv_dumper_2378;
    csv_file_dump cstatus_csv_dumper_2378;
    df_fifo_monitor fifo_monitor_2378;
    df_fifo_intf fifo_intf_2379(clock,reset);
    assign fifo_intf_2379.rd_en = AESL_inst_myproject.layer3_out_1026_U.if_read & AESL_inst_myproject.layer3_out_1026_U.if_empty_n;
    assign fifo_intf_2379.wr_en = AESL_inst_myproject.layer3_out_1026_U.if_write & AESL_inst_myproject.layer3_out_1026_U.if_full_n;
    assign fifo_intf_2379.fifo_rd_block = 0;
    assign fifo_intf_2379.fifo_wr_block = 0;
    assign fifo_intf_2379.finish = finish;
    csv_file_dump fifo_csv_dumper_2379;
    csv_file_dump cstatus_csv_dumper_2379;
    df_fifo_monitor fifo_monitor_2379;
    df_fifo_intf fifo_intf_2380(clock,reset);
    assign fifo_intf_2380.rd_en = AESL_inst_myproject.layer3_out_1027_U.if_read & AESL_inst_myproject.layer3_out_1027_U.if_empty_n;
    assign fifo_intf_2380.wr_en = AESL_inst_myproject.layer3_out_1027_U.if_write & AESL_inst_myproject.layer3_out_1027_U.if_full_n;
    assign fifo_intf_2380.fifo_rd_block = 0;
    assign fifo_intf_2380.fifo_wr_block = 0;
    assign fifo_intf_2380.finish = finish;
    csv_file_dump fifo_csv_dumper_2380;
    csv_file_dump cstatus_csv_dumper_2380;
    df_fifo_monitor fifo_monitor_2380;
    df_fifo_intf fifo_intf_2381(clock,reset);
    assign fifo_intf_2381.rd_en = AESL_inst_myproject.layer3_out_1028_U.if_read & AESL_inst_myproject.layer3_out_1028_U.if_empty_n;
    assign fifo_intf_2381.wr_en = AESL_inst_myproject.layer3_out_1028_U.if_write & AESL_inst_myproject.layer3_out_1028_U.if_full_n;
    assign fifo_intf_2381.fifo_rd_block = 0;
    assign fifo_intf_2381.fifo_wr_block = 0;
    assign fifo_intf_2381.finish = finish;
    csv_file_dump fifo_csv_dumper_2381;
    csv_file_dump cstatus_csv_dumper_2381;
    df_fifo_monitor fifo_monitor_2381;
    df_fifo_intf fifo_intf_2382(clock,reset);
    assign fifo_intf_2382.rd_en = AESL_inst_myproject.layer3_out_1029_U.if_read & AESL_inst_myproject.layer3_out_1029_U.if_empty_n;
    assign fifo_intf_2382.wr_en = AESL_inst_myproject.layer3_out_1029_U.if_write & AESL_inst_myproject.layer3_out_1029_U.if_full_n;
    assign fifo_intf_2382.fifo_rd_block = 0;
    assign fifo_intf_2382.fifo_wr_block = 0;
    assign fifo_intf_2382.finish = finish;
    csv_file_dump fifo_csv_dumper_2382;
    csv_file_dump cstatus_csv_dumper_2382;
    df_fifo_monitor fifo_monitor_2382;
    df_fifo_intf fifo_intf_2383(clock,reset);
    assign fifo_intf_2383.rd_en = AESL_inst_myproject.layer3_out_1030_U.if_read & AESL_inst_myproject.layer3_out_1030_U.if_empty_n;
    assign fifo_intf_2383.wr_en = AESL_inst_myproject.layer3_out_1030_U.if_write & AESL_inst_myproject.layer3_out_1030_U.if_full_n;
    assign fifo_intf_2383.fifo_rd_block = 0;
    assign fifo_intf_2383.fifo_wr_block = 0;
    assign fifo_intf_2383.finish = finish;
    csv_file_dump fifo_csv_dumper_2383;
    csv_file_dump cstatus_csv_dumper_2383;
    df_fifo_monitor fifo_monitor_2383;
    df_fifo_intf fifo_intf_2384(clock,reset);
    assign fifo_intf_2384.rd_en = AESL_inst_myproject.layer3_out_1031_U.if_read & AESL_inst_myproject.layer3_out_1031_U.if_empty_n;
    assign fifo_intf_2384.wr_en = AESL_inst_myproject.layer3_out_1031_U.if_write & AESL_inst_myproject.layer3_out_1031_U.if_full_n;
    assign fifo_intf_2384.fifo_rd_block = 0;
    assign fifo_intf_2384.fifo_wr_block = 0;
    assign fifo_intf_2384.finish = finish;
    csv_file_dump fifo_csv_dumper_2384;
    csv_file_dump cstatus_csv_dumper_2384;
    df_fifo_monitor fifo_monitor_2384;
    df_fifo_intf fifo_intf_2385(clock,reset);
    assign fifo_intf_2385.rd_en = AESL_inst_myproject.layer3_out_1032_U.if_read & AESL_inst_myproject.layer3_out_1032_U.if_empty_n;
    assign fifo_intf_2385.wr_en = AESL_inst_myproject.layer3_out_1032_U.if_write & AESL_inst_myproject.layer3_out_1032_U.if_full_n;
    assign fifo_intf_2385.fifo_rd_block = 0;
    assign fifo_intf_2385.fifo_wr_block = 0;
    assign fifo_intf_2385.finish = finish;
    csv_file_dump fifo_csv_dumper_2385;
    csv_file_dump cstatus_csv_dumper_2385;
    df_fifo_monitor fifo_monitor_2385;
    df_fifo_intf fifo_intf_2386(clock,reset);
    assign fifo_intf_2386.rd_en = AESL_inst_myproject.layer3_out_1033_U.if_read & AESL_inst_myproject.layer3_out_1033_U.if_empty_n;
    assign fifo_intf_2386.wr_en = AESL_inst_myproject.layer3_out_1033_U.if_write & AESL_inst_myproject.layer3_out_1033_U.if_full_n;
    assign fifo_intf_2386.fifo_rd_block = 0;
    assign fifo_intf_2386.fifo_wr_block = 0;
    assign fifo_intf_2386.finish = finish;
    csv_file_dump fifo_csv_dumper_2386;
    csv_file_dump cstatus_csv_dumper_2386;
    df_fifo_monitor fifo_monitor_2386;
    df_fifo_intf fifo_intf_2387(clock,reset);
    assign fifo_intf_2387.rd_en = AESL_inst_myproject.layer3_out_1034_U.if_read & AESL_inst_myproject.layer3_out_1034_U.if_empty_n;
    assign fifo_intf_2387.wr_en = AESL_inst_myproject.layer3_out_1034_U.if_write & AESL_inst_myproject.layer3_out_1034_U.if_full_n;
    assign fifo_intf_2387.fifo_rd_block = 0;
    assign fifo_intf_2387.fifo_wr_block = 0;
    assign fifo_intf_2387.finish = finish;
    csv_file_dump fifo_csv_dumper_2387;
    csv_file_dump cstatus_csv_dumper_2387;
    df_fifo_monitor fifo_monitor_2387;
    df_fifo_intf fifo_intf_2388(clock,reset);
    assign fifo_intf_2388.rd_en = AESL_inst_myproject.layer3_out_1035_U.if_read & AESL_inst_myproject.layer3_out_1035_U.if_empty_n;
    assign fifo_intf_2388.wr_en = AESL_inst_myproject.layer3_out_1035_U.if_write & AESL_inst_myproject.layer3_out_1035_U.if_full_n;
    assign fifo_intf_2388.fifo_rd_block = 0;
    assign fifo_intf_2388.fifo_wr_block = 0;
    assign fifo_intf_2388.finish = finish;
    csv_file_dump fifo_csv_dumper_2388;
    csv_file_dump cstatus_csv_dumper_2388;
    df_fifo_monitor fifo_monitor_2388;
    df_fifo_intf fifo_intf_2389(clock,reset);
    assign fifo_intf_2389.rd_en = AESL_inst_myproject.layer3_out_1036_U.if_read & AESL_inst_myproject.layer3_out_1036_U.if_empty_n;
    assign fifo_intf_2389.wr_en = AESL_inst_myproject.layer3_out_1036_U.if_write & AESL_inst_myproject.layer3_out_1036_U.if_full_n;
    assign fifo_intf_2389.fifo_rd_block = 0;
    assign fifo_intf_2389.fifo_wr_block = 0;
    assign fifo_intf_2389.finish = finish;
    csv_file_dump fifo_csv_dumper_2389;
    csv_file_dump cstatus_csv_dumper_2389;
    df_fifo_monitor fifo_monitor_2389;
    df_fifo_intf fifo_intf_2390(clock,reset);
    assign fifo_intf_2390.rd_en = AESL_inst_myproject.layer3_out_1037_U.if_read & AESL_inst_myproject.layer3_out_1037_U.if_empty_n;
    assign fifo_intf_2390.wr_en = AESL_inst_myproject.layer3_out_1037_U.if_write & AESL_inst_myproject.layer3_out_1037_U.if_full_n;
    assign fifo_intf_2390.fifo_rd_block = 0;
    assign fifo_intf_2390.fifo_wr_block = 0;
    assign fifo_intf_2390.finish = finish;
    csv_file_dump fifo_csv_dumper_2390;
    csv_file_dump cstatus_csv_dumper_2390;
    df_fifo_monitor fifo_monitor_2390;
    df_fifo_intf fifo_intf_2391(clock,reset);
    assign fifo_intf_2391.rd_en = AESL_inst_myproject.layer3_out_1038_U.if_read & AESL_inst_myproject.layer3_out_1038_U.if_empty_n;
    assign fifo_intf_2391.wr_en = AESL_inst_myproject.layer3_out_1038_U.if_write & AESL_inst_myproject.layer3_out_1038_U.if_full_n;
    assign fifo_intf_2391.fifo_rd_block = 0;
    assign fifo_intf_2391.fifo_wr_block = 0;
    assign fifo_intf_2391.finish = finish;
    csv_file_dump fifo_csv_dumper_2391;
    csv_file_dump cstatus_csv_dumper_2391;
    df_fifo_monitor fifo_monitor_2391;
    df_fifo_intf fifo_intf_2392(clock,reset);
    assign fifo_intf_2392.rd_en = AESL_inst_myproject.layer3_out_1039_U.if_read & AESL_inst_myproject.layer3_out_1039_U.if_empty_n;
    assign fifo_intf_2392.wr_en = AESL_inst_myproject.layer3_out_1039_U.if_write & AESL_inst_myproject.layer3_out_1039_U.if_full_n;
    assign fifo_intf_2392.fifo_rd_block = 0;
    assign fifo_intf_2392.fifo_wr_block = 0;
    assign fifo_intf_2392.finish = finish;
    csv_file_dump fifo_csv_dumper_2392;
    csv_file_dump cstatus_csv_dumper_2392;
    df_fifo_monitor fifo_monitor_2392;
    df_fifo_intf fifo_intf_2393(clock,reset);
    assign fifo_intf_2393.rd_en = AESL_inst_myproject.layer3_out_1040_U.if_read & AESL_inst_myproject.layer3_out_1040_U.if_empty_n;
    assign fifo_intf_2393.wr_en = AESL_inst_myproject.layer3_out_1040_U.if_write & AESL_inst_myproject.layer3_out_1040_U.if_full_n;
    assign fifo_intf_2393.fifo_rd_block = 0;
    assign fifo_intf_2393.fifo_wr_block = 0;
    assign fifo_intf_2393.finish = finish;
    csv_file_dump fifo_csv_dumper_2393;
    csv_file_dump cstatus_csv_dumper_2393;
    df_fifo_monitor fifo_monitor_2393;
    df_fifo_intf fifo_intf_2394(clock,reset);
    assign fifo_intf_2394.rd_en = AESL_inst_myproject.layer3_out_1041_U.if_read & AESL_inst_myproject.layer3_out_1041_U.if_empty_n;
    assign fifo_intf_2394.wr_en = AESL_inst_myproject.layer3_out_1041_U.if_write & AESL_inst_myproject.layer3_out_1041_U.if_full_n;
    assign fifo_intf_2394.fifo_rd_block = 0;
    assign fifo_intf_2394.fifo_wr_block = 0;
    assign fifo_intf_2394.finish = finish;
    csv_file_dump fifo_csv_dumper_2394;
    csv_file_dump cstatus_csv_dumper_2394;
    df_fifo_monitor fifo_monitor_2394;
    df_fifo_intf fifo_intf_2395(clock,reset);
    assign fifo_intf_2395.rd_en = AESL_inst_myproject.layer3_out_1042_U.if_read & AESL_inst_myproject.layer3_out_1042_U.if_empty_n;
    assign fifo_intf_2395.wr_en = AESL_inst_myproject.layer3_out_1042_U.if_write & AESL_inst_myproject.layer3_out_1042_U.if_full_n;
    assign fifo_intf_2395.fifo_rd_block = 0;
    assign fifo_intf_2395.fifo_wr_block = 0;
    assign fifo_intf_2395.finish = finish;
    csv_file_dump fifo_csv_dumper_2395;
    csv_file_dump cstatus_csv_dumper_2395;
    df_fifo_monitor fifo_monitor_2395;
    df_fifo_intf fifo_intf_2396(clock,reset);
    assign fifo_intf_2396.rd_en = AESL_inst_myproject.layer3_out_1043_U.if_read & AESL_inst_myproject.layer3_out_1043_U.if_empty_n;
    assign fifo_intf_2396.wr_en = AESL_inst_myproject.layer3_out_1043_U.if_write & AESL_inst_myproject.layer3_out_1043_U.if_full_n;
    assign fifo_intf_2396.fifo_rd_block = 0;
    assign fifo_intf_2396.fifo_wr_block = 0;
    assign fifo_intf_2396.finish = finish;
    csv_file_dump fifo_csv_dumper_2396;
    csv_file_dump cstatus_csv_dumper_2396;
    df_fifo_monitor fifo_monitor_2396;
    df_fifo_intf fifo_intf_2397(clock,reset);
    assign fifo_intf_2397.rd_en = AESL_inst_myproject.layer3_out_1044_U.if_read & AESL_inst_myproject.layer3_out_1044_U.if_empty_n;
    assign fifo_intf_2397.wr_en = AESL_inst_myproject.layer3_out_1044_U.if_write & AESL_inst_myproject.layer3_out_1044_U.if_full_n;
    assign fifo_intf_2397.fifo_rd_block = 0;
    assign fifo_intf_2397.fifo_wr_block = 0;
    assign fifo_intf_2397.finish = finish;
    csv_file_dump fifo_csv_dumper_2397;
    csv_file_dump cstatus_csv_dumper_2397;
    df_fifo_monitor fifo_monitor_2397;
    df_fifo_intf fifo_intf_2398(clock,reset);
    assign fifo_intf_2398.rd_en = AESL_inst_myproject.layer3_out_1045_U.if_read & AESL_inst_myproject.layer3_out_1045_U.if_empty_n;
    assign fifo_intf_2398.wr_en = AESL_inst_myproject.layer3_out_1045_U.if_write & AESL_inst_myproject.layer3_out_1045_U.if_full_n;
    assign fifo_intf_2398.fifo_rd_block = 0;
    assign fifo_intf_2398.fifo_wr_block = 0;
    assign fifo_intf_2398.finish = finish;
    csv_file_dump fifo_csv_dumper_2398;
    csv_file_dump cstatus_csv_dumper_2398;
    df_fifo_monitor fifo_monitor_2398;
    df_fifo_intf fifo_intf_2399(clock,reset);
    assign fifo_intf_2399.rd_en = AESL_inst_myproject.layer3_out_1046_U.if_read & AESL_inst_myproject.layer3_out_1046_U.if_empty_n;
    assign fifo_intf_2399.wr_en = AESL_inst_myproject.layer3_out_1046_U.if_write & AESL_inst_myproject.layer3_out_1046_U.if_full_n;
    assign fifo_intf_2399.fifo_rd_block = 0;
    assign fifo_intf_2399.fifo_wr_block = 0;
    assign fifo_intf_2399.finish = finish;
    csv_file_dump fifo_csv_dumper_2399;
    csv_file_dump cstatus_csv_dumper_2399;
    df_fifo_monitor fifo_monitor_2399;
    df_fifo_intf fifo_intf_2400(clock,reset);
    assign fifo_intf_2400.rd_en = AESL_inst_myproject.layer3_out_1047_U.if_read & AESL_inst_myproject.layer3_out_1047_U.if_empty_n;
    assign fifo_intf_2400.wr_en = AESL_inst_myproject.layer3_out_1047_U.if_write & AESL_inst_myproject.layer3_out_1047_U.if_full_n;
    assign fifo_intf_2400.fifo_rd_block = 0;
    assign fifo_intf_2400.fifo_wr_block = 0;
    assign fifo_intf_2400.finish = finish;
    csv_file_dump fifo_csv_dumper_2400;
    csv_file_dump cstatus_csv_dumper_2400;
    df_fifo_monitor fifo_monitor_2400;
    df_fifo_intf fifo_intf_2401(clock,reset);
    assign fifo_intf_2401.rd_en = AESL_inst_myproject.layer3_out_1048_U.if_read & AESL_inst_myproject.layer3_out_1048_U.if_empty_n;
    assign fifo_intf_2401.wr_en = AESL_inst_myproject.layer3_out_1048_U.if_write & AESL_inst_myproject.layer3_out_1048_U.if_full_n;
    assign fifo_intf_2401.fifo_rd_block = 0;
    assign fifo_intf_2401.fifo_wr_block = 0;
    assign fifo_intf_2401.finish = finish;
    csv_file_dump fifo_csv_dumper_2401;
    csv_file_dump cstatus_csv_dumper_2401;
    df_fifo_monitor fifo_monitor_2401;
    df_fifo_intf fifo_intf_2402(clock,reset);
    assign fifo_intf_2402.rd_en = AESL_inst_myproject.layer3_out_1049_U.if_read & AESL_inst_myproject.layer3_out_1049_U.if_empty_n;
    assign fifo_intf_2402.wr_en = AESL_inst_myproject.layer3_out_1049_U.if_write & AESL_inst_myproject.layer3_out_1049_U.if_full_n;
    assign fifo_intf_2402.fifo_rd_block = 0;
    assign fifo_intf_2402.fifo_wr_block = 0;
    assign fifo_intf_2402.finish = finish;
    csv_file_dump fifo_csv_dumper_2402;
    csv_file_dump cstatus_csv_dumper_2402;
    df_fifo_monitor fifo_monitor_2402;
    df_fifo_intf fifo_intf_2403(clock,reset);
    assign fifo_intf_2403.rd_en = AESL_inst_myproject.layer3_out_1050_U.if_read & AESL_inst_myproject.layer3_out_1050_U.if_empty_n;
    assign fifo_intf_2403.wr_en = AESL_inst_myproject.layer3_out_1050_U.if_write & AESL_inst_myproject.layer3_out_1050_U.if_full_n;
    assign fifo_intf_2403.fifo_rd_block = 0;
    assign fifo_intf_2403.fifo_wr_block = 0;
    assign fifo_intf_2403.finish = finish;
    csv_file_dump fifo_csv_dumper_2403;
    csv_file_dump cstatus_csv_dumper_2403;
    df_fifo_monitor fifo_monitor_2403;
    df_fifo_intf fifo_intf_2404(clock,reset);
    assign fifo_intf_2404.rd_en = AESL_inst_myproject.layer3_out_1051_U.if_read & AESL_inst_myproject.layer3_out_1051_U.if_empty_n;
    assign fifo_intf_2404.wr_en = AESL_inst_myproject.layer3_out_1051_U.if_write & AESL_inst_myproject.layer3_out_1051_U.if_full_n;
    assign fifo_intf_2404.fifo_rd_block = 0;
    assign fifo_intf_2404.fifo_wr_block = 0;
    assign fifo_intf_2404.finish = finish;
    csv_file_dump fifo_csv_dumper_2404;
    csv_file_dump cstatus_csv_dumper_2404;
    df_fifo_monitor fifo_monitor_2404;
    df_fifo_intf fifo_intf_2405(clock,reset);
    assign fifo_intf_2405.rd_en = AESL_inst_myproject.layer3_out_1052_U.if_read & AESL_inst_myproject.layer3_out_1052_U.if_empty_n;
    assign fifo_intf_2405.wr_en = AESL_inst_myproject.layer3_out_1052_U.if_write & AESL_inst_myproject.layer3_out_1052_U.if_full_n;
    assign fifo_intf_2405.fifo_rd_block = 0;
    assign fifo_intf_2405.fifo_wr_block = 0;
    assign fifo_intf_2405.finish = finish;
    csv_file_dump fifo_csv_dumper_2405;
    csv_file_dump cstatus_csv_dumper_2405;
    df_fifo_monitor fifo_monitor_2405;
    df_fifo_intf fifo_intf_2406(clock,reset);
    assign fifo_intf_2406.rd_en = AESL_inst_myproject.layer3_out_1053_U.if_read & AESL_inst_myproject.layer3_out_1053_U.if_empty_n;
    assign fifo_intf_2406.wr_en = AESL_inst_myproject.layer3_out_1053_U.if_write & AESL_inst_myproject.layer3_out_1053_U.if_full_n;
    assign fifo_intf_2406.fifo_rd_block = 0;
    assign fifo_intf_2406.fifo_wr_block = 0;
    assign fifo_intf_2406.finish = finish;
    csv_file_dump fifo_csv_dumper_2406;
    csv_file_dump cstatus_csv_dumper_2406;
    df_fifo_monitor fifo_monitor_2406;
    df_fifo_intf fifo_intf_2407(clock,reset);
    assign fifo_intf_2407.rd_en = AESL_inst_myproject.layer3_out_1054_U.if_read & AESL_inst_myproject.layer3_out_1054_U.if_empty_n;
    assign fifo_intf_2407.wr_en = AESL_inst_myproject.layer3_out_1054_U.if_write & AESL_inst_myproject.layer3_out_1054_U.if_full_n;
    assign fifo_intf_2407.fifo_rd_block = 0;
    assign fifo_intf_2407.fifo_wr_block = 0;
    assign fifo_intf_2407.finish = finish;
    csv_file_dump fifo_csv_dumper_2407;
    csv_file_dump cstatus_csv_dumper_2407;
    df_fifo_monitor fifo_monitor_2407;
    df_fifo_intf fifo_intf_2408(clock,reset);
    assign fifo_intf_2408.rd_en = AESL_inst_myproject.layer3_out_1055_U.if_read & AESL_inst_myproject.layer3_out_1055_U.if_empty_n;
    assign fifo_intf_2408.wr_en = AESL_inst_myproject.layer3_out_1055_U.if_write & AESL_inst_myproject.layer3_out_1055_U.if_full_n;
    assign fifo_intf_2408.fifo_rd_block = 0;
    assign fifo_intf_2408.fifo_wr_block = 0;
    assign fifo_intf_2408.finish = finish;
    csv_file_dump fifo_csv_dumper_2408;
    csv_file_dump cstatus_csv_dumper_2408;
    df_fifo_monitor fifo_monitor_2408;
    df_fifo_intf fifo_intf_2409(clock,reset);
    assign fifo_intf_2409.rd_en = AESL_inst_myproject.layer3_out_1056_U.if_read & AESL_inst_myproject.layer3_out_1056_U.if_empty_n;
    assign fifo_intf_2409.wr_en = AESL_inst_myproject.layer3_out_1056_U.if_write & AESL_inst_myproject.layer3_out_1056_U.if_full_n;
    assign fifo_intf_2409.fifo_rd_block = 0;
    assign fifo_intf_2409.fifo_wr_block = 0;
    assign fifo_intf_2409.finish = finish;
    csv_file_dump fifo_csv_dumper_2409;
    csv_file_dump cstatus_csv_dumper_2409;
    df_fifo_monitor fifo_monitor_2409;
    df_fifo_intf fifo_intf_2410(clock,reset);
    assign fifo_intf_2410.rd_en = AESL_inst_myproject.layer3_out_1057_U.if_read & AESL_inst_myproject.layer3_out_1057_U.if_empty_n;
    assign fifo_intf_2410.wr_en = AESL_inst_myproject.layer3_out_1057_U.if_write & AESL_inst_myproject.layer3_out_1057_U.if_full_n;
    assign fifo_intf_2410.fifo_rd_block = 0;
    assign fifo_intf_2410.fifo_wr_block = 0;
    assign fifo_intf_2410.finish = finish;
    csv_file_dump fifo_csv_dumper_2410;
    csv_file_dump cstatus_csv_dumper_2410;
    df_fifo_monitor fifo_monitor_2410;
    df_fifo_intf fifo_intf_2411(clock,reset);
    assign fifo_intf_2411.rd_en = AESL_inst_myproject.layer3_out_1058_U.if_read & AESL_inst_myproject.layer3_out_1058_U.if_empty_n;
    assign fifo_intf_2411.wr_en = AESL_inst_myproject.layer3_out_1058_U.if_write & AESL_inst_myproject.layer3_out_1058_U.if_full_n;
    assign fifo_intf_2411.fifo_rd_block = 0;
    assign fifo_intf_2411.fifo_wr_block = 0;
    assign fifo_intf_2411.finish = finish;
    csv_file_dump fifo_csv_dumper_2411;
    csv_file_dump cstatus_csv_dumper_2411;
    df_fifo_monitor fifo_monitor_2411;
    df_fifo_intf fifo_intf_2412(clock,reset);
    assign fifo_intf_2412.rd_en = AESL_inst_myproject.layer3_out_1059_U.if_read & AESL_inst_myproject.layer3_out_1059_U.if_empty_n;
    assign fifo_intf_2412.wr_en = AESL_inst_myproject.layer3_out_1059_U.if_write & AESL_inst_myproject.layer3_out_1059_U.if_full_n;
    assign fifo_intf_2412.fifo_rd_block = 0;
    assign fifo_intf_2412.fifo_wr_block = 0;
    assign fifo_intf_2412.finish = finish;
    csv_file_dump fifo_csv_dumper_2412;
    csv_file_dump cstatus_csv_dumper_2412;
    df_fifo_monitor fifo_monitor_2412;
    df_fifo_intf fifo_intf_2413(clock,reset);
    assign fifo_intf_2413.rd_en = AESL_inst_myproject.layer3_out_1060_U.if_read & AESL_inst_myproject.layer3_out_1060_U.if_empty_n;
    assign fifo_intf_2413.wr_en = AESL_inst_myproject.layer3_out_1060_U.if_write & AESL_inst_myproject.layer3_out_1060_U.if_full_n;
    assign fifo_intf_2413.fifo_rd_block = 0;
    assign fifo_intf_2413.fifo_wr_block = 0;
    assign fifo_intf_2413.finish = finish;
    csv_file_dump fifo_csv_dumper_2413;
    csv_file_dump cstatus_csv_dumper_2413;
    df_fifo_monitor fifo_monitor_2413;
    df_fifo_intf fifo_intf_2414(clock,reset);
    assign fifo_intf_2414.rd_en = AESL_inst_myproject.layer3_out_1061_U.if_read & AESL_inst_myproject.layer3_out_1061_U.if_empty_n;
    assign fifo_intf_2414.wr_en = AESL_inst_myproject.layer3_out_1061_U.if_write & AESL_inst_myproject.layer3_out_1061_U.if_full_n;
    assign fifo_intf_2414.fifo_rd_block = 0;
    assign fifo_intf_2414.fifo_wr_block = 0;
    assign fifo_intf_2414.finish = finish;
    csv_file_dump fifo_csv_dumper_2414;
    csv_file_dump cstatus_csv_dumper_2414;
    df_fifo_monitor fifo_monitor_2414;
    df_fifo_intf fifo_intf_2415(clock,reset);
    assign fifo_intf_2415.rd_en = AESL_inst_myproject.layer3_out_1062_U.if_read & AESL_inst_myproject.layer3_out_1062_U.if_empty_n;
    assign fifo_intf_2415.wr_en = AESL_inst_myproject.layer3_out_1062_U.if_write & AESL_inst_myproject.layer3_out_1062_U.if_full_n;
    assign fifo_intf_2415.fifo_rd_block = 0;
    assign fifo_intf_2415.fifo_wr_block = 0;
    assign fifo_intf_2415.finish = finish;
    csv_file_dump fifo_csv_dumper_2415;
    csv_file_dump cstatus_csv_dumper_2415;
    df_fifo_monitor fifo_monitor_2415;
    df_fifo_intf fifo_intf_2416(clock,reset);
    assign fifo_intf_2416.rd_en = AESL_inst_myproject.layer3_out_1063_U.if_read & AESL_inst_myproject.layer3_out_1063_U.if_empty_n;
    assign fifo_intf_2416.wr_en = AESL_inst_myproject.layer3_out_1063_U.if_write & AESL_inst_myproject.layer3_out_1063_U.if_full_n;
    assign fifo_intf_2416.fifo_rd_block = 0;
    assign fifo_intf_2416.fifo_wr_block = 0;
    assign fifo_intf_2416.finish = finish;
    csv_file_dump fifo_csv_dumper_2416;
    csv_file_dump cstatus_csv_dumper_2416;
    df_fifo_monitor fifo_monitor_2416;
    df_fifo_intf fifo_intf_2417(clock,reset);
    assign fifo_intf_2417.rd_en = AESL_inst_myproject.layer3_out_1064_U.if_read & AESL_inst_myproject.layer3_out_1064_U.if_empty_n;
    assign fifo_intf_2417.wr_en = AESL_inst_myproject.layer3_out_1064_U.if_write & AESL_inst_myproject.layer3_out_1064_U.if_full_n;
    assign fifo_intf_2417.fifo_rd_block = 0;
    assign fifo_intf_2417.fifo_wr_block = 0;
    assign fifo_intf_2417.finish = finish;
    csv_file_dump fifo_csv_dumper_2417;
    csv_file_dump cstatus_csv_dumper_2417;
    df_fifo_monitor fifo_monitor_2417;
    df_fifo_intf fifo_intf_2418(clock,reset);
    assign fifo_intf_2418.rd_en = AESL_inst_myproject.layer3_out_1065_U.if_read & AESL_inst_myproject.layer3_out_1065_U.if_empty_n;
    assign fifo_intf_2418.wr_en = AESL_inst_myproject.layer3_out_1065_U.if_write & AESL_inst_myproject.layer3_out_1065_U.if_full_n;
    assign fifo_intf_2418.fifo_rd_block = 0;
    assign fifo_intf_2418.fifo_wr_block = 0;
    assign fifo_intf_2418.finish = finish;
    csv_file_dump fifo_csv_dumper_2418;
    csv_file_dump cstatus_csv_dumper_2418;
    df_fifo_monitor fifo_monitor_2418;
    df_fifo_intf fifo_intf_2419(clock,reset);
    assign fifo_intf_2419.rd_en = AESL_inst_myproject.layer3_out_1066_U.if_read & AESL_inst_myproject.layer3_out_1066_U.if_empty_n;
    assign fifo_intf_2419.wr_en = AESL_inst_myproject.layer3_out_1066_U.if_write & AESL_inst_myproject.layer3_out_1066_U.if_full_n;
    assign fifo_intf_2419.fifo_rd_block = 0;
    assign fifo_intf_2419.fifo_wr_block = 0;
    assign fifo_intf_2419.finish = finish;
    csv_file_dump fifo_csv_dumper_2419;
    csv_file_dump cstatus_csv_dumper_2419;
    df_fifo_monitor fifo_monitor_2419;
    df_fifo_intf fifo_intf_2420(clock,reset);
    assign fifo_intf_2420.rd_en = AESL_inst_myproject.layer3_out_1067_U.if_read & AESL_inst_myproject.layer3_out_1067_U.if_empty_n;
    assign fifo_intf_2420.wr_en = AESL_inst_myproject.layer3_out_1067_U.if_write & AESL_inst_myproject.layer3_out_1067_U.if_full_n;
    assign fifo_intf_2420.fifo_rd_block = 0;
    assign fifo_intf_2420.fifo_wr_block = 0;
    assign fifo_intf_2420.finish = finish;
    csv_file_dump fifo_csv_dumper_2420;
    csv_file_dump cstatus_csv_dumper_2420;
    df_fifo_monitor fifo_monitor_2420;
    df_fifo_intf fifo_intf_2421(clock,reset);
    assign fifo_intf_2421.rd_en = AESL_inst_myproject.layer3_out_1068_U.if_read & AESL_inst_myproject.layer3_out_1068_U.if_empty_n;
    assign fifo_intf_2421.wr_en = AESL_inst_myproject.layer3_out_1068_U.if_write & AESL_inst_myproject.layer3_out_1068_U.if_full_n;
    assign fifo_intf_2421.fifo_rd_block = 0;
    assign fifo_intf_2421.fifo_wr_block = 0;
    assign fifo_intf_2421.finish = finish;
    csv_file_dump fifo_csv_dumper_2421;
    csv_file_dump cstatus_csv_dumper_2421;
    df_fifo_monitor fifo_monitor_2421;
    df_fifo_intf fifo_intf_2422(clock,reset);
    assign fifo_intf_2422.rd_en = AESL_inst_myproject.layer3_out_1069_U.if_read & AESL_inst_myproject.layer3_out_1069_U.if_empty_n;
    assign fifo_intf_2422.wr_en = AESL_inst_myproject.layer3_out_1069_U.if_write & AESL_inst_myproject.layer3_out_1069_U.if_full_n;
    assign fifo_intf_2422.fifo_rd_block = 0;
    assign fifo_intf_2422.fifo_wr_block = 0;
    assign fifo_intf_2422.finish = finish;
    csv_file_dump fifo_csv_dumper_2422;
    csv_file_dump cstatus_csv_dumper_2422;
    df_fifo_monitor fifo_monitor_2422;
    df_fifo_intf fifo_intf_2423(clock,reset);
    assign fifo_intf_2423.rd_en = AESL_inst_myproject.layer3_out_1070_U.if_read & AESL_inst_myproject.layer3_out_1070_U.if_empty_n;
    assign fifo_intf_2423.wr_en = AESL_inst_myproject.layer3_out_1070_U.if_write & AESL_inst_myproject.layer3_out_1070_U.if_full_n;
    assign fifo_intf_2423.fifo_rd_block = 0;
    assign fifo_intf_2423.fifo_wr_block = 0;
    assign fifo_intf_2423.finish = finish;
    csv_file_dump fifo_csv_dumper_2423;
    csv_file_dump cstatus_csv_dumper_2423;
    df_fifo_monitor fifo_monitor_2423;
    df_fifo_intf fifo_intf_2424(clock,reset);
    assign fifo_intf_2424.rd_en = AESL_inst_myproject.layer3_out_1071_U.if_read & AESL_inst_myproject.layer3_out_1071_U.if_empty_n;
    assign fifo_intf_2424.wr_en = AESL_inst_myproject.layer3_out_1071_U.if_write & AESL_inst_myproject.layer3_out_1071_U.if_full_n;
    assign fifo_intf_2424.fifo_rd_block = 0;
    assign fifo_intf_2424.fifo_wr_block = 0;
    assign fifo_intf_2424.finish = finish;
    csv_file_dump fifo_csv_dumper_2424;
    csv_file_dump cstatus_csv_dumper_2424;
    df_fifo_monitor fifo_monitor_2424;
    df_fifo_intf fifo_intf_2425(clock,reset);
    assign fifo_intf_2425.rd_en = AESL_inst_myproject.layer3_out_1072_U.if_read & AESL_inst_myproject.layer3_out_1072_U.if_empty_n;
    assign fifo_intf_2425.wr_en = AESL_inst_myproject.layer3_out_1072_U.if_write & AESL_inst_myproject.layer3_out_1072_U.if_full_n;
    assign fifo_intf_2425.fifo_rd_block = 0;
    assign fifo_intf_2425.fifo_wr_block = 0;
    assign fifo_intf_2425.finish = finish;
    csv_file_dump fifo_csv_dumper_2425;
    csv_file_dump cstatus_csv_dumper_2425;
    df_fifo_monitor fifo_monitor_2425;
    df_fifo_intf fifo_intf_2426(clock,reset);
    assign fifo_intf_2426.rd_en = AESL_inst_myproject.layer3_out_1073_U.if_read & AESL_inst_myproject.layer3_out_1073_U.if_empty_n;
    assign fifo_intf_2426.wr_en = AESL_inst_myproject.layer3_out_1073_U.if_write & AESL_inst_myproject.layer3_out_1073_U.if_full_n;
    assign fifo_intf_2426.fifo_rd_block = 0;
    assign fifo_intf_2426.fifo_wr_block = 0;
    assign fifo_intf_2426.finish = finish;
    csv_file_dump fifo_csv_dumper_2426;
    csv_file_dump cstatus_csv_dumper_2426;
    df_fifo_monitor fifo_monitor_2426;
    df_fifo_intf fifo_intf_2427(clock,reset);
    assign fifo_intf_2427.rd_en = AESL_inst_myproject.layer3_out_1074_U.if_read & AESL_inst_myproject.layer3_out_1074_U.if_empty_n;
    assign fifo_intf_2427.wr_en = AESL_inst_myproject.layer3_out_1074_U.if_write & AESL_inst_myproject.layer3_out_1074_U.if_full_n;
    assign fifo_intf_2427.fifo_rd_block = 0;
    assign fifo_intf_2427.fifo_wr_block = 0;
    assign fifo_intf_2427.finish = finish;
    csv_file_dump fifo_csv_dumper_2427;
    csv_file_dump cstatus_csv_dumper_2427;
    df_fifo_monitor fifo_monitor_2427;
    df_fifo_intf fifo_intf_2428(clock,reset);
    assign fifo_intf_2428.rd_en = AESL_inst_myproject.layer3_out_1075_U.if_read & AESL_inst_myproject.layer3_out_1075_U.if_empty_n;
    assign fifo_intf_2428.wr_en = AESL_inst_myproject.layer3_out_1075_U.if_write & AESL_inst_myproject.layer3_out_1075_U.if_full_n;
    assign fifo_intf_2428.fifo_rd_block = 0;
    assign fifo_intf_2428.fifo_wr_block = 0;
    assign fifo_intf_2428.finish = finish;
    csv_file_dump fifo_csv_dumper_2428;
    csv_file_dump cstatus_csv_dumper_2428;
    df_fifo_monitor fifo_monitor_2428;
    df_fifo_intf fifo_intf_2429(clock,reset);
    assign fifo_intf_2429.rd_en = AESL_inst_myproject.layer3_out_1076_U.if_read & AESL_inst_myproject.layer3_out_1076_U.if_empty_n;
    assign fifo_intf_2429.wr_en = AESL_inst_myproject.layer3_out_1076_U.if_write & AESL_inst_myproject.layer3_out_1076_U.if_full_n;
    assign fifo_intf_2429.fifo_rd_block = 0;
    assign fifo_intf_2429.fifo_wr_block = 0;
    assign fifo_intf_2429.finish = finish;
    csv_file_dump fifo_csv_dumper_2429;
    csv_file_dump cstatus_csv_dumper_2429;
    df_fifo_monitor fifo_monitor_2429;
    df_fifo_intf fifo_intf_2430(clock,reset);
    assign fifo_intf_2430.rd_en = AESL_inst_myproject.layer3_out_1077_U.if_read & AESL_inst_myproject.layer3_out_1077_U.if_empty_n;
    assign fifo_intf_2430.wr_en = AESL_inst_myproject.layer3_out_1077_U.if_write & AESL_inst_myproject.layer3_out_1077_U.if_full_n;
    assign fifo_intf_2430.fifo_rd_block = 0;
    assign fifo_intf_2430.fifo_wr_block = 0;
    assign fifo_intf_2430.finish = finish;
    csv_file_dump fifo_csv_dumper_2430;
    csv_file_dump cstatus_csv_dumper_2430;
    df_fifo_monitor fifo_monitor_2430;
    df_fifo_intf fifo_intf_2431(clock,reset);
    assign fifo_intf_2431.rd_en = AESL_inst_myproject.layer3_out_1078_U.if_read & AESL_inst_myproject.layer3_out_1078_U.if_empty_n;
    assign fifo_intf_2431.wr_en = AESL_inst_myproject.layer3_out_1078_U.if_write & AESL_inst_myproject.layer3_out_1078_U.if_full_n;
    assign fifo_intf_2431.fifo_rd_block = 0;
    assign fifo_intf_2431.fifo_wr_block = 0;
    assign fifo_intf_2431.finish = finish;
    csv_file_dump fifo_csv_dumper_2431;
    csv_file_dump cstatus_csv_dumper_2431;
    df_fifo_monitor fifo_monitor_2431;
    df_fifo_intf fifo_intf_2432(clock,reset);
    assign fifo_intf_2432.rd_en = AESL_inst_myproject.layer3_out_1079_U.if_read & AESL_inst_myproject.layer3_out_1079_U.if_empty_n;
    assign fifo_intf_2432.wr_en = AESL_inst_myproject.layer3_out_1079_U.if_write & AESL_inst_myproject.layer3_out_1079_U.if_full_n;
    assign fifo_intf_2432.fifo_rd_block = 0;
    assign fifo_intf_2432.fifo_wr_block = 0;
    assign fifo_intf_2432.finish = finish;
    csv_file_dump fifo_csv_dumper_2432;
    csv_file_dump cstatus_csv_dumper_2432;
    df_fifo_monitor fifo_monitor_2432;
    df_fifo_intf fifo_intf_2433(clock,reset);
    assign fifo_intf_2433.rd_en = AESL_inst_myproject.layer3_out_1080_U.if_read & AESL_inst_myproject.layer3_out_1080_U.if_empty_n;
    assign fifo_intf_2433.wr_en = AESL_inst_myproject.layer3_out_1080_U.if_write & AESL_inst_myproject.layer3_out_1080_U.if_full_n;
    assign fifo_intf_2433.fifo_rd_block = 0;
    assign fifo_intf_2433.fifo_wr_block = 0;
    assign fifo_intf_2433.finish = finish;
    csv_file_dump fifo_csv_dumper_2433;
    csv_file_dump cstatus_csv_dumper_2433;
    df_fifo_monitor fifo_monitor_2433;
    df_fifo_intf fifo_intf_2434(clock,reset);
    assign fifo_intf_2434.rd_en = AESL_inst_myproject.layer3_out_1081_U.if_read & AESL_inst_myproject.layer3_out_1081_U.if_empty_n;
    assign fifo_intf_2434.wr_en = AESL_inst_myproject.layer3_out_1081_U.if_write & AESL_inst_myproject.layer3_out_1081_U.if_full_n;
    assign fifo_intf_2434.fifo_rd_block = 0;
    assign fifo_intf_2434.fifo_wr_block = 0;
    assign fifo_intf_2434.finish = finish;
    csv_file_dump fifo_csv_dumper_2434;
    csv_file_dump cstatus_csv_dumper_2434;
    df_fifo_monitor fifo_monitor_2434;
    df_fifo_intf fifo_intf_2435(clock,reset);
    assign fifo_intf_2435.rd_en = AESL_inst_myproject.layer3_out_1082_U.if_read & AESL_inst_myproject.layer3_out_1082_U.if_empty_n;
    assign fifo_intf_2435.wr_en = AESL_inst_myproject.layer3_out_1082_U.if_write & AESL_inst_myproject.layer3_out_1082_U.if_full_n;
    assign fifo_intf_2435.fifo_rd_block = 0;
    assign fifo_intf_2435.fifo_wr_block = 0;
    assign fifo_intf_2435.finish = finish;
    csv_file_dump fifo_csv_dumper_2435;
    csv_file_dump cstatus_csv_dumper_2435;
    df_fifo_monitor fifo_monitor_2435;
    df_fifo_intf fifo_intf_2436(clock,reset);
    assign fifo_intf_2436.rd_en = AESL_inst_myproject.layer3_out_1083_U.if_read & AESL_inst_myproject.layer3_out_1083_U.if_empty_n;
    assign fifo_intf_2436.wr_en = AESL_inst_myproject.layer3_out_1083_U.if_write & AESL_inst_myproject.layer3_out_1083_U.if_full_n;
    assign fifo_intf_2436.fifo_rd_block = 0;
    assign fifo_intf_2436.fifo_wr_block = 0;
    assign fifo_intf_2436.finish = finish;
    csv_file_dump fifo_csv_dumper_2436;
    csv_file_dump cstatus_csv_dumper_2436;
    df_fifo_monitor fifo_monitor_2436;
    df_fifo_intf fifo_intf_2437(clock,reset);
    assign fifo_intf_2437.rd_en = AESL_inst_myproject.layer3_out_1084_U.if_read & AESL_inst_myproject.layer3_out_1084_U.if_empty_n;
    assign fifo_intf_2437.wr_en = AESL_inst_myproject.layer3_out_1084_U.if_write & AESL_inst_myproject.layer3_out_1084_U.if_full_n;
    assign fifo_intf_2437.fifo_rd_block = 0;
    assign fifo_intf_2437.fifo_wr_block = 0;
    assign fifo_intf_2437.finish = finish;
    csv_file_dump fifo_csv_dumper_2437;
    csv_file_dump cstatus_csv_dumper_2437;
    df_fifo_monitor fifo_monitor_2437;
    df_fifo_intf fifo_intf_2438(clock,reset);
    assign fifo_intf_2438.rd_en = AESL_inst_myproject.layer3_out_1085_U.if_read & AESL_inst_myproject.layer3_out_1085_U.if_empty_n;
    assign fifo_intf_2438.wr_en = AESL_inst_myproject.layer3_out_1085_U.if_write & AESL_inst_myproject.layer3_out_1085_U.if_full_n;
    assign fifo_intf_2438.fifo_rd_block = 0;
    assign fifo_intf_2438.fifo_wr_block = 0;
    assign fifo_intf_2438.finish = finish;
    csv_file_dump fifo_csv_dumper_2438;
    csv_file_dump cstatus_csv_dumper_2438;
    df_fifo_monitor fifo_monitor_2438;
    df_fifo_intf fifo_intf_2439(clock,reset);
    assign fifo_intf_2439.rd_en = AESL_inst_myproject.layer3_out_1086_U.if_read & AESL_inst_myproject.layer3_out_1086_U.if_empty_n;
    assign fifo_intf_2439.wr_en = AESL_inst_myproject.layer3_out_1086_U.if_write & AESL_inst_myproject.layer3_out_1086_U.if_full_n;
    assign fifo_intf_2439.fifo_rd_block = 0;
    assign fifo_intf_2439.fifo_wr_block = 0;
    assign fifo_intf_2439.finish = finish;
    csv_file_dump fifo_csv_dumper_2439;
    csv_file_dump cstatus_csv_dumper_2439;
    df_fifo_monitor fifo_monitor_2439;
    df_fifo_intf fifo_intf_2440(clock,reset);
    assign fifo_intf_2440.rd_en = AESL_inst_myproject.layer3_out_1087_U.if_read & AESL_inst_myproject.layer3_out_1087_U.if_empty_n;
    assign fifo_intf_2440.wr_en = AESL_inst_myproject.layer3_out_1087_U.if_write & AESL_inst_myproject.layer3_out_1087_U.if_full_n;
    assign fifo_intf_2440.fifo_rd_block = 0;
    assign fifo_intf_2440.fifo_wr_block = 0;
    assign fifo_intf_2440.finish = finish;
    csv_file_dump fifo_csv_dumper_2440;
    csv_file_dump cstatus_csv_dumper_2440;
    df_fifo_monitor fifo_monitor_2440;
    df_fifo_intf fifo_intf_2441(clock,reset);
    assign fifo_intf_2441.rd_en = AESL_inst_myproject.layer3_out_1088_U.if_read & AESL_inst_myproject.layer3_out_1088_U.if_empty_n;
    assign fifo_intf_2441.wr_en = AESL_inst_myproject.layer3_out_1088_U.if_write & AESL_inst_myproject.layer3_out_1088_U.if_full_n;
    assign fifo_intf_2441.fifo_rd_block = 0;
    assign fifo_intf_2441.fifo_wr_block = 0;
    assign fifo_intf_2441.finish = finish;
    csv_file_dump fifo_csv_dumper_2441;
    csv_file_dump cstatus_csv_dumper_2441;
    df_fifo_monitor fifo_monitor_2441;
    df_fifo_intf fifo_intf_2442(clock,reset);
    assign fifo_intf_2442.rd_en = AESL_inst_myproject.layer3_out_1089_U.if_read & AESL_inst_myproject.layer3_out_1089_U.if_empty_n;
    assign fifo_intf_2442.wr_en = AESL_inst_myproject.layer3_out_1089_U.if_write & AESL_inst_myproject.layer3_out_1089_U.if_full_n;
    assign fifo_intf_2442.fifo_rd_block = 0;
    assign fifo_intf_2442.fifo_wr_block = 0;
    assign fifo_intf_2442.finish = finish;
    csv_file_dump fifo_csv_dumper_2442;
    csv_file_dump cstatus_csv_dumper_2442;
    df_fifo_monitor fifo_monitor_2442;
    df_fifo_intf fifo_intf_2443(clock,reset);
    assign fifo_intf_2443.rd_en = AESL_inst_myproject.layer3_out_1090_U.if_read & AESL_inst_myproject.layer3_out_1090_U.if_empty_n;
    assign fifo_intf_2443.wr_en = AESL_inst_myproject.layer3_out_1090_U.if_write & AESL_inst_myproject.layer3_out_1090_U.if_full_n;
    assign fifo_intf_2443.fifo_rd_block = 0;
    assign fifo_intf_2443.fifo_wr_block = 0;
    assign fifo_intf_2443.finish = finish;
    csv_file_dump fifo_csv_dumper_2443;
    csv_file_dump cstatus_csv_dumper_2443;
    df_fifo_monitor fifo_monitor_2443;
    df_fifo_intf fifo_intf_2444(clock,reset);
    assign fifo_intf_2444.rd_en = AESL_inst_myproject.layer3_out_1091_U.if_read & AESL_inst_myproject.layer3_out_1091_U.if_empty_n;
    assign fifo_intf_2444.wr_en = AESL_inst_myproject.layer3_out_1091_U.if_write & AESL_inst_myproject.layer3_out_1091_U.if_full_n;
    assign fifo_intf_2444.fifo_rd_block = 0;
    assign fifo_intf_2444.fifo_wr_block = 0;
    assign fifo_intf_2444.finish = finish;
    csv_file_dump fifo_csv_dumper_2444;
    csv_file_dump cstatus_csv_dumper_2444;
    df_fifo_monitor fifo_monitor_2444;
    df_fifo_intf fifo_intf_2445(clock,reset);
    assign fifo_intf_2445.rd_en = AESL_inst_myproject.layer3_out_1092_U.if_read & AESL_inst_myproject.layer3_out_1092_U.if_empty_n;
    assign fifo_intf_2445.wr_en = AESL_inst_myproject.layer3_out_1092_U.if_write & AESL_inst_myproject.layer3_out_1092_U.if_full_n;
    assign fifo_intf_2445.fifo_rd_block = 0;
    assign fifo_intf_2445.fifo_wr_block = 0;
    assign fifo_intf_2445.finish = finish;
    csv_file_dump fifo_csv_dumper_2445;
    csv_file_dump cstatus_csv_dumper_2445;
    df_fifo_monitor fifo_monitor_2445;
    df_fifo_intf fifo_intf_2446(clock,reset);
    assign fifo_intf_2446.rd_en = AESL_inst_myproject.layer3_out_1093_U.if_read & AESL_inst_myproject.layer3_out_1093_U.if_empty_n;
    assign fifo_intf_2446.wr_en = AESL_inst_myproject.layer3_out_1093_U.if_write & AESL_inst_myproject.layer3_out_1093_U.if_full_n;
    assign fifo_intf_2446.fifo_rd_block = 0;
    assign fifo_intf_2446.fifo_wr_block = 0;
    assign fifo_intf_2446.finish = finish;
    csv_file_dump fifo_csv_dumper_2446;
    csv_file_dump cstatus_csv_dumper_2446;
    df_fifo_monitor fifo_monitor_2446;
    df_fifo_intf fifo_intf_2447(clock,reset);
    assign fifo_intf_2447.rd_en = AESL_inst_myproject.layer3_out_1094_U.if_read & AESL_inst_myproject.layer3_out_1094_U.if_empty_n;
    assign fifo_intf_2447.wr_en = AESL_inst_myproject.layer3_out_1094_U.if_write & AESL_inst_myproject.layer3_out_1094_U.if_full_n;
    assign fifo_intf_2447.fifo_rd_block = 0;
    assign fifo_intf_2447.fifo_wr_block = 0;
    assign fifo_intf_2447.finish = finish;
    csv_file_dump fifo_csv_dumper_2447;
    csv_file_dump cstatus_csv_dumper_2447;
    df_fifo_monitor fifo_monitor_2447;
    df_fifo_intf fifo_intf_2448(clock,reset);
    assign fifo_intf_2448.rd_en = AESL_inst_myproject.layer3_out_1095_U.if_read & AESL_inst_myproject.layer3_out_1095_U.if_empty_n;
    assign fifo_intf_2448.wr_en = AESL_inst_myproject.layer3_out_1095_U.if_write & AESL_inst_myproject.layer3_out_1095_U.if_full_n;
    assign fifo_intf_2448.fifo_rd_block = 0;
    assign fifo_intf_2448.fifo_wr_block = 0;
    assign fifo_intf_2448.finish = finish;
    csv_file_dump fifo_csv_dumper_2448;
    csv_file_dump cstatus_csv_dumper_2448;
    df_fifo_monitor fifo_monitor_2448;
    df_fifo_intf fifo_intf_2449(clock,reset);
    assign fifo_intf_2449.rd_en = AESL_inst_myproject.layer3_out_1096_U.if_read & AESL_inst_myproject.layer3_out_1096_U.if_empty_n;
    assign fifo_intf_2449.wr_en = AESL_inst_myproject.layer3_out_1096_U.if_write & AESL_inst_myproject.layer3_out_1096_U.if_full_n;
    assign fifo_intf_2449.fifo_rd_block = 0;
    assign fifo_intf_2449.fifo_wr_block = 0;
    assign fifo_intf_2449.finish = finish;
    csv_file_dump fifo_csv_dumper_2449;
    csv_file_dump cstatus_csv_dumper_2449;
    df_fifo_monitor fifo_monitor_2449;
    df_fifo_intf fifo_intf_2450(clock,reset);
    assign fifo_intf_2450.rd_en = AESL_inst_myproject.layer3_out_1097_U.if_read & AESL_inst_myproject.layer3_out_1097_U.if_empty_n;
    assign fifo_intf_2450.wr_en = AESL_inst_myproject.layer3_out_1097_U.if_write & AESL_inst_myproject.layer3_out_1097_U.if_full_n;
    assign fifo_intf_2450.fifo_rd_block = 0;
    assign fifo_intf_2450.fifo_wr_block = 0;
    assign fifo_intf_2450.finish = finish;
    csv_file_dump fifo_csv_dumper_2450;
    csv_file_dump cstatus_csv_dumper_2450;
    df_fifo_monitor fifo_monitor_2450;
    df_fifo_intf fifo_intf_2451(clock,reset);
    assign fifo_intf_2451.rd_en = AESL_inst_myproject.layer3_out_1098_U.if_read & AESL_inst_myproject.layer3_out_1098_U.if_empty_n;
    assign fifo_intf_2451.wr_en = AESL_inst_myproject.layer3_out_1098_U.if_write & AESL_inst_myproject.layer3_out_1098_U.if_full_n;
    assign fifo_intf_2451.fifo_rd_block = 0;
    assign fifo_intf_2451.fifo_wr_block = 0;
    assign fifo_intf_2451.finish = finish;
    csv_file_dump fifo_csv_dumper_2451;
    csv_file_dump cstatus_csv_dumper_2451;
    df_fifo_monitor fifo_monitor_2451;
    df_fifo_intf fifo_intf_2452(clock,reset);
    assign fifo_intf_2452.rd_en = AESL_inst_myproject.layer3_out_1099_U.if_read & AESL_inst_myproject.layer3_out_1099_U.if_empty_n;
    assign fifo_intf_2452.wr_en = AESL_inst_myproject.layer3_out_1099_U.if_write & AESL_inst_myproject.layer3_out_1099_U.if_full_n;
    assign fifo_intf_2452.fifo_rd_block = 0;
    assign fifo_intf_2452.fifo_wr_block = 0;
    assign fifo_intf_2452.finish = finish;
    csv_file_dump fifo_csv_dumper_2452;
    csv_file_dump cstatus_csv_dumper_2452;
    df_fifo_monitor fifo_monitor_2452;
    df_fifo_intf fifo_intf_2453(clock,reset);
    assign fifo_intf_2453.rd_en = AESL_inst_myproject.layer3_out_1100_U.if_read & AESL_inst_myproject.layer3_out_1100_U.if_empty_n;
    assign fifo_intf_2453.wr_en = AESL_inst_myproject.layer3_out_1100_U.if_write & AESL_inst_myproject.layer3_out_1100_U.if_full_n;
    assign fifo_intf_2453.fifo_rd_block = 0;
    assign fifo_intf_2453.fifo_wr_block = 0;
    assign fifo_intf_2453.finish = finish;
    csv_file_dump fifo_csv_dumper_2453;
    csv_file_dump cstatus_csv_dumper_2453;
    df_fifo_monitor fifo_monitor_2453;
    df_fifo_intf fifo_intf_2454(clock,reset);
    assign fifo_intf_2454.rd_en = AESL_inst_myproject.layer3_out_1101_U.if_read & AESL_inst_myproject.layer3_out_1101_U.if_empty_n;
    assign fifo_intf_2454.wr_en = AESL_inst_myproject.layer3_out_1101_U.if_write & AESL_inst_myproject.layer3_out_1101_U.if_full_n;
    assign fifo_intf_2454.fifo_rd_block = 0;
    assign fifo_intf_2454.fifo_wr_block = 0;
    assign fifo_intf_2454.finish = finish;
    csv_file_dump fifo_csv_dumper_2454;
    csv_file_dump cstatus_csv_dumper_2454;
    df_fifo_monitor fifo_monitor_2454;
    df_fifo_intf fifo_intf_2455(clock,reset);
    assign fifo_intf_2455.rd_en = AESL_inst_myproject.layer3_out_1102_U.if_read & AESL_inst_myproject.layer3_out_1102_U.if_empty_n;
    assign fifo_intf_2455.wr_en = AESL_inst_myproject.layer3_out_1102_U.if_write & AESL_inst_myproject.layer3_out_1102_U.if_full_n;
    assign fifo_intf_2455.fifo_rd_block = 0;
    assign fifo_intf_2455.fifo_wr_block = 0;
    assign fifo_intf_2455.finish = finish;
    csv_file_dump fifo_csv_dumper_2455;
    csv_file_dump cstatus_csv_dumper_2455;
    df_fifo_monitor fifo_monitor_2455;
    df_fifo_intf fifo_intf_2456(clock,reset);
    assign fifo_intf_2456.rd_en = AESL_inst_myproject.layer3_out_1103_U.if_read & AESL_inst_myproject.layer3_out_1103_U.if_empty_n;
    assign fifo_intf_2456.wr_en = AESL_inst_myproject.layer3_out_1103_U.if_write & AESL_inst_myproject.layer3_out_1103_U.if_full_n;
    assign fifo_intf_2456.fifo_rd_block = 0;
    assign fifo_intf_2456.fifo_wr_block = 0;
    assign fifo_intf_2456.finish = finish;
    csv_file_dump fifo_csv_dumper_2456;
    csv_file_dump cstatus_csv_dumper_2456;
    df_fifo_monitor fifo_monitor_2456;
    df_fifo_intf fifo_intf_2457(clock,reset);
    assign fifo_intf_2457.rd_en = AESL_inst_myproject.layer3_out_1104_U.if_read & AESL_inst_myproject.layer3_out_1104_U.if_empty_n;
    assign fifo_intf_2457.wr_en = AESL_inst_myproject.layer3_out_1104_U.if_write & AESL_inst_myproject.layer3_out_1104_U.if_full_n;
    assign fifo_intf_2457.fifo_rd_block = 0;
    assign fifo_intf_2457.fifo_wr_block = 0;
    assign fifo_intf_2457.finish = finish;
    csv_file_dump fifo_csv_dumper_2457;
    csv_file_dump cstatus_csv_dumper_2457;
    df_fifo_monitor fifo_monitor_2457;
    df_fifo_intf fifo_intf_2458(clock,reset);
    assign fifo_intf_2458.rd_en = AESL_inst_myproject.layer3_out_1105_U.if_read & AESL_inst_myproject.layer3_out_1105_U.if_empty_n;
    assign fifo_intf_2458.wr_en = AESL_inst_myproject.layer3_out_1105_U.if_write & AESL_inst_myproject.layer3_out_1105_U.if_full_n;
    assign fifo_intf_2458.fifo_rd_block = 0;
    assign fifo_intf_2458.fifo_wr_block = 0;
    assign fifo_intf_2458.finish = finish;
    csv_file_dump fifo_csv_dumper_2458;
    csv_file_dump cstatus_csv_dumper_2458;
    df_fifo_monitor fifo_monitor_2458;
    df_fifo_intf fifo_intf_2459(clock,reset);
    assign fifo_intf_2459.rd_en = AESL_inst_myproject.layer3_out_1106_U.if_read & AESL_inst_myproject.layer3_out_1106_U.if_empty_n;
    assign fifo_intf_2459.wr_en = AESL_inst_myproject.layer3_out_1106_U.if_write & AESL_inst_myproject.layer3_out_1106_U.if_full_n;
    assign fifo_intf_2459.fifo_rd_block = 0;
    assign fifo_intf_2459.fifo_wr_block = 0;
    assign fifo_intf_2459.finish = finish;
    csv_file_dump fifo_csv_dumper_2459;
    csv_file_dump cstatus_csv_dumper_2459;
    df_fifo_monitor fifo_monitor_2459;
    df_fifo_intf fifo_intf_2460(clock,reset);
    assign fifo_intf_2460.rd_en = AESL_inst_myproject.layer3_out_1107_U.if_read & AESL_inst_myproject.layer3_out_1107_U.if_empty_n;
    assign fifo_intf_2460.wr_en = AESL_inst_myproject.layer3_out_1107_U.if_write & AESL_inst_myproject.layer3_out_1107_U.if_full_n;
    assign fifo_intf_2460.fifo_rd_block = 0;
    assign fifo_intf_2460.fifo_wr_block = 0;
    assign fifo_intf_2460.finish = finish;
    csv_file_dump fifo_csv_dumper_2460;
    csv_file_dump cstatus_csv_dumper_2460;
    df_fifo_monitor fifo_monitor_2460;
    df_fifo_intf fifo_intf_2461(clock,reset);
    assign fifo_intf_2461.rd_en = AESL_inst_myproject.layer3_out_1108_U.if_read & AESL_inst_myproject.layer3_out_1108_U.if_empty_n;
    assign fifo_intf_2461.wr_en = AESL_inst_myproject.layer3_out_1108_U.if_write & AESL_inst_myproject.layer3_out_1108_U.if_full_n;
    assign fifo_intf_2461.fifo_rd_block = 0;
    assign fifo_intf_2461.fifo_wr_block = 0;
    assign fifo_intf_2461.finish = finish;
    csv_file_dump fifo_csv_dumper_2461;
    csv_file_dump cstatus_csv_dumper_2461;
    df_fifo_monitor fifo_monitor_2461;
    df_fifo_intf fifo_intf_2462(clock,reset);
    assign fifo_intf_2462.rd_en = AESL_inst_myproject.layer3_out_1109_U.if_read & AESL_inst_myproject.layer3_out_1109_U.if_empty_n;
    assign fifo_intf_2462.wr_en = AESL_inst_myproject.layer3_out_1109_U.if_write & AESL_inst_myproject.layer3_out_1109_U.if_full_n;
    assign fifo_intf_2462.fifo_rd_block = 0;
    assign fifo_intf_2462.fifo_wr_block = 0;
    assign fifo_intf_2462.finish = finish;
    csv_file_dump fifo_csv_dumper_2462;
    csv_file_dump cstatus_csv_dumper_2462;
    df_fifo_monitor fifo_monitor_2462;
    df_fifo_intf fifo_intf_2463(clock,reset);
    assign fifo_intf_2463.rd_en = AESL_inst_myproject.layer3_out_1110_U.if_read & AESL_inst_myproject.layer3_out_1110_U.if_empty_n;
    assign fifo_intf_2463.wr_en = AESL_inst_myproject.layer3_out_1110_U.if_write & AESL_inst_myproject.layer3_out_1110_U.if_full_n;
    assign fifo_intf_2463.fifo_rd_block = 0;
    assign fifo_intf_2463.fifo_wr_block = 0;
    assign fifo_intf_2463.finish = finish;
    csv_file_dump fifo_csv_dumper_2463;
    csv_file_dump cstatus_csv_dumper_2463;
    df_fifo_monitor fifo_monitor_2463;
    df_fifo_intf fifo_intf_2464(clock,reset);
    assign fifo_intf_2464.rd_en = AESL_inst_myproject.layer3_out_1111_U.if_read & AESL_inst_myproject.layer3_out_1111_U.if_empty_n;
    assign fifo_intf_2464.wr_en = AESL_inst_myproject.layer3_out_1111_U.if_write & AESL_inst_myproject.layer3_out_1111_U.if_full_n;
    assign fifo_intf_2464.fifo_rd_block = 0;
    assign fifo_intf_2464.fifo_wr_block = 0;
    assign fifo_intf_2464.finish = finish;
    csv_file_dump fifo_csv_dumper_2464;
    csv_file_dump cstatus_csv_dumper_2464;
    df_fifo_monitor fifo_monitor_2464;
    df_fifo_intf fifo_intf_2465(clock,reset);
    assign fifo_intf_2465.rd_en = AESL_inst_myproject.layer3_out_1112_U.if_read & AESL_inst_myproject.layer3_out_1112_U.if_empty_n;
    assign fifo_intf_2465.wr_en = AESL_inst_myproject.layer3_out_1112_U.if_write & AESL_inst_myproject.layer3_out_1112_U.if_full_n;
    assign fifo_intf_2465.fifo_rd_block = 0;
    assign fifo_intf_2465.fifo_wr_block = 0;
    assign fifo_intf_2465.finish = finish;
    csv_file_dump fifo_csv_dumper_2465;
    csv_file_dump cstatus_csv_dumper_2465;
    df_fifo_monitor fifo_monitor_2465;
    df_fifo_intf fifo_intf_2466(clock,reset);
    assign fifo_intf_2466.rd_en = AESL_inst_myproject.layer3_out_1113_U.if_read & AESL_inst_myproject.layer3_out_1113_U.if_empty_n;
    assign fifo_intf_2466.wr_en = AESL_inst_myproject.layer3_out_1113_U.if_write & AESL_inst_myproject.layer3_out_1113_U.if_full_n;
    assign fifo_intf_2466.fifo_rd_block = 0;
    assign fifo_intf_2466.fifo_wr_block = 0;
    assign fifo_intf_2466.finish = finish;
    csv_file_dump fifo_csv_dumper_2466;
    csv_file_dump cstatus_csv_dumper_2466;
    df_fifo_monitor fifo_monitor_2466;
    df_fifo_intf fifo_intf_2467(clock,reset);
    assign fifo_intf_2467.rd_en = AESL_inst_myproject.layer3_out_1114_U.if_read & AESL_inst_myproject.layer3_out_1114_U.if_empty_n;
    assign fifo_intf_2467.wr_en = AESL_inst_myproject.layer3_out_1114_U.if_write & AESL_inst_myproject.layer3_out_1114_U.if_full_n;
    assign fifo_intf_2467.fifo_rd_block = 0;
    assign fifo_intf_2467.fifo_wr_block = 0;
    assign fifo_intf_2467.finish = finish;
    csv_file_dump fifo_csv_dumper_2467;
    csv_file_dump cstatus_csv_dumper_2467;
    df_fifo_monitor fifo_monitor_2467;
    df_fifo_intf fifo_intf_2468(clock,reset);
    assign fifo_intf_2468.rd_en = AESL_inst_myproject.layer3_out_1115_U.if_read & AESL_inst_myproject.layer3_out_1115_U.if_empty_n;
    assign fifo_intf_2468.wr_en = AESL_inst_myproject.layer3_out_1115_U.if_write & AESL_inst_myproject.layer3_out_1115_U.if_full_n;
    assign fifo_intf_2468.fifo_rd_block = 0;
    assign fifo_intf_2468.fifo_wr_block = 0;
    assign fifo_intf_2468.finish = finish;
    csv_file_dump fifo_csv_dumper_2468;
    csv_file_dump cstatus_csv_dumper_2468;
    df_fifo_monitor fifo_monitor_2468;
    df_fifo_intf fifo_intf_2469(clock,reset);
    assign fifo_intf_2469.rd_en = AESL_inst_myproject.layer3_out_1116_U.if_read & AESL_inst_myproject.layer3_out_1116_U.if_empty_n;
    assign fifo_intf_2469.wr_en = AESL_inst_myproject.layer3_out_1116_U.if_write & AESL_inst_myproject.layer3_out_1116_U.if_full_n;
    assign fifo_intf_2469.fifo_rd_block = 0;
    assign fifo_intf_2469.fifo_wr_block = 0;
    assign fifo_intf_2469.finish = finish;
    csv_file_dump fifo_csv_dumper_2469;
    csv_file_dump cstatus_csv_dumper_2469;
    df_fifo_monitor fifo_monitor_2469;
    df_fifo_intf fifo_intf_2470(clock,reset);
    assign fifo_intf_2470.rd_en = AESL_inst_myproject.layer3_out_1117_U.if_read & AESL_inst_myproject.layer3_out_1117_U.if_empty_n;
    assign fifo_intf_2470.wr_en = AESL_inst_myproject.layer3_out_1117_U.if_write & AESL_inst_myproject.layer3_out_1117_U.if_full_n;
    assign fifo_intf_2470.fifo_rd_block = 0;
    assign fifo_intf_2470.fifo_wr_block = 0;
    assign fifo_intf_2470.finish = finish;
    csv_file_dump fifo_csv_dumper_2470;
    csv_file_dump cstatus_csv_dumper_2470;
    df_fifo_monitor fifo_monitor_2470;
    df_fifo_intf fifo_intf_2471(clock,reset);
    assign fifo_intf_2471.rd_en = AESL_inst_myproject.layer3_out_1118_U.if_read & AESL_inst_myproject.layer3_out_1118_U.if_empty_n;
    assign fifo_intf_2471.wr_en = AESL_inst_myproject.layer3_out_1118_U.if_write & AESL_inst_myproject.layer3_out_1118_U.if_full_n;
    assign fifo_intf_2471.fifo_rd_block = 0;
    assign fifo_intf_2471.fifo_wr_block = 0;
    assign fifo_intf_2471.finish = finish;
    csv_file_dump fifo_csv_dumper_2471;
    csv_file_dump cstatus_csv_dumper_2471;
    df_fifo_monitor fifo_monitor_2471;
    df_fifo_intf fifo_intf_2472(clock,reset);
    assign fifo_intf_2472.rd_en = AESL_inst_myproject.layer3_out_1119_U.if_read & AESL_inst_myproject.layer3_out_1119_U.if_empty_n;
    assign fifo_intf_2472.wr_en = AESL_inst_myproject.layer3_out_1119_U.if_write & AESL_inst_myproject.layer3_out_1119_U.if_full_n;
    assign fifo_intf_2472.fifo_rd_block = 0;
    assign fifo_intf_2472.fifo_wr_block = 0;
    assign fifo_intf_2472.finish = finish;
    csv_file_dump fifo_csv_dumper_2472;
    csv_file_dump cstatus_csv_dumper_2472;
    df_fifo_monitor fifo_monitor_2472;
    df_fifo_intf fifo_intf_2473(clock,reset);
    assign fifo_intf_2473.rd_en = AESL_inst_myproject.layer3_out_1120_U.if_read & AESL_inst_myproject.layer3_out_1120_U.if_empty_n;
    assign fifo_intf_2473.wr_en = AESL_inst_myproject.layer3_out_1120_U.if_write & AESL_inst_myproject.layer3_out_1120_U.if_full_n;
    assign fifo_intf_2473.fifo_rd_block = 0;
    assign fifo_intf_2473.fifo_wr_block = 0;
    assign fifo_intf_2473.finish = finish;
    csv_file_dump fifo_csv_dumper_2473;
    csv_file_dump cstatus_csv_dumper_2473;
    df_fifo_monitor fifo_monitor_2473;
    df_fifo_intf fifo_intf_2474(clock,reset);
    assign fifo_intf_2474.rd_en = AESL_inst_myproject.layer3_out_1121_U.if_read & AESL_inst_myproject.layer3_out_1121_U.if_empty_n;
    assign fifo_intf_2474.wr_en = AESL_inst_myproject.layer3_out_1121_U.if_write & AESL_inst_myproject.layer3_out_1121_U.if_full_n;
    assign fifo_intf_2474.fifo_rd_block = 0;
    assign fifo_intf_2474.fifo_wr_block = 0;
    assign fifo_intf_2474.finish = finish;
    csv_file_dump fifo_csv_dumper_2474;
    csv_file_dump cstatus_csv_dumper_2474;
    df_fifo_monitor fifo_monitor_2474;
    df_fifo_intf fifo_intf_2475(clock,reset);
    assign fifo_intf_2475.rd_en = AESL_inst_myproject.layer3_out_1122_U.if_read & AESL_inst_myproject.layer3_out_1122_U.if_empty_n;
    assign fifo_intf_2475.wr_en = AESL_inst_myproject.layer3_out_1122_U.if_write & AESL_inst_myproject.layer3_out_1122_U.if_full_n;
    assign fifo_intf_2475.fifo_rd_block = 0;
    assign fifo_intf_2475.fifo_wr_block = 0;
    assign fifo_intf_2475.finish = finish;
    csv_file_dump fifo_csv_dumper_2475;
    csv_file_dump cstatus_csv_dumper_2475;
    df_fifo_monitor fifo_monitor_2475;
    df_fifo_intf fifo_intf_2476(clock,reset);
    assign fifo_intf_2476.rd_en = AESL_inst_myproject.layer3_out_1123_U.if_read & AESL_inst_myproject.layer3_out_1123_U.if_empty_n;
    assign fifo_intf_2476.wr_en = AESL_inst_myproject.layer3_out_1123_U.if_write & AESL_inst_myproject.layer3_out_1123_U.if_full_n;
    assign fifo_intf_2476.fifo_rd_block = 0;
    assign fifo_intf_2476.fifo_wr_block = 0;
    assign fifo_intf_2476.finish = finish;
    csv_file_dump fifo_csv_dumper_2476;
    csv_file_dump cstatus_csv_dumper_2476;
    df_fifo_monitor fifo_monitor_2476;
    df_fifo_intf fifo_intf_2477(clock,reset);
    assign fifo_intf_2477.rd_en = AESL_inst_myproject.layer3_out_1124_U.if_read & AESL_inst_myproject.layer3_out_1124_U.if_empty_n;
    assign fifo_intf_2477.wr_en = AESL_inst_myproject.layer3_out_1124_U.if_write & AESL_inst_myproject.layer3_out_1124_U.if_full_n;
    assign fifo_intf_2477.fifo_rd_block = 0;
    assign fifo_intf_2477.fifo_wr_block = 0;
    assign fifo_intf_2477.finish = finish;
    csv_file_dump fifo_csv_dumper_2477;
    csv_file_dump cstatus_csv_dumper_2477;
    df_fifo_monitor fifo_monitor_2477;
    df_fifo_intf fifo_intf_2478(clock,reset);
    assign fifo_intf_2478.rd_en = AESL_inst_myproject.layer3_out_1125_U.if_read & AESL_inst_myproject.layer3_out_1125_U.if_empty_n;
    assign fifo_intf_2478.wr_en = AESL_inst_myproject.layer3_out_1125_U.if_write & AESL_inst_myproject.layer3_out_1125_U.if_full_n;
    assign fifo_intf_2478.fifo_rd_block = 0;
    assign fifo_intf_2478.fifo_wr_block = 0;
    assign fifo_intf_2478.finish = finish;
    csv_file_dump fifo_csv_dumper_2478;
    csv_file_dump cstatus_csv_dumper_2478;
    df_fifo_monitor fifo_monitor_2478;
    df_fifo_intf fifo_intf_2479(clock,reset);
    assign fifo_intf_2479.rd_en = AESL_inst_myproject.layer3_out_1126_U.if_read & AESL_inst_myproject.layer3_out_1126_U.if_empty_n;
    assign fifo_intf_2479.wr_en = AESL_inst_myproject.layer3_out_1126_U.if_write & AESL_inst_myproject.layer3_out_1126_U.if_full_n;
    assign fifo_intf_2479.fifo_rd_block = 0;
    assign fifo_intf_2479.fifo_wr_block = 0;
    assign fifo_intf_2479.finish = finish;
    csv_file_dump fifo_csv_dumper_2479;
    csv_file_dump cstatus_csv_dumper_2479;
    df_fifo_monitor fifo_monitor_2479;
    df_fifo_intf fifo_intf_2480(clock,reset);
    assign fifo_intf_2480.rd_en = AESL_inst_myproject.layer3_out_1127_U.if_read & AESL_inst_myproject.layer3_out_1127_U.if_empty_n;
    assign fifo_intf_2480.wr_en = AESL_inst_myproject.layer3_out_1127_U.if_write & AESL_inst_myproject.layer3_out_1127_U.if_full_n;
    assign fifo_intf_2480.fifo_rd_block = 0;
    assign fifo_intf_2480.fifo_wr_block = 0;
    assign fifo_intf_2480.finish = finish;
    csv_file_dump fifo_csv_dumper_2480;
    csv_file_dump cstatus_csv_dumper_2480;
    df_fifo_monitor fifo_monitor_2480;
    df_fifo_intf fifo_intf_2481(clock,reset);
    assign fifo_intf_2481.rd_en = AESL_inst_myproject.layer3_out_1128_U.if_read & AESL_inst_myproject.layer3_out_1128_U.if_empty_n;
    assign fifo_intf_2481.wr_en = AESL_inst_myproject.layer3_out_1128_U.if_write & AESL_inst_myproject.layer3_out_1128_U.if_full_n;
    assign fifo_intf_2481.fifo_rd_block = 0;
    assign fifo_intf_2481.fifo_wr_block = 0;
    assign fifo_intf_2481.finish = finish;
    csv_file_dump fifo_csv_dumper_2481;
    csv_file_dump cstatus_csv_dumper_2481;
    df_fifo_monitor fifo_monitor_2481;
    df_fifo_intf fifo_intf_2482(clock,reset);
    assign fifo_intf_2482.rd_en = AESL_inst_myproject.layer3_out_1129_U.if_read & AESL_inst_myproject.layer3_out_1129_U.if_empty_n;
    assign fifo_intf_2482.wr_en = AESL_inst_myproject.layer3_out_1129_U.if_write & AESL_inst_myproject.layer3_out_1129_U.if_full_n;
    assign fifo_intf_2482.fifo_rd_block = 0;
    assign fifo_intf_2482.fifo_wr_block = 0;
    assign fifo_intf_2482.finish = finish;
    csv_file_dump fifo_csv_dumper_2482;
    csv_file_dump cstatus_csv_dumper_2482;
    df_fifo_monitor fifo_monitor_2482;
    df_fifo_intf fifo_intf_2483(clock,reset);
    assign fifo_intf_2483.rd_en = AESL_inst_myproject.layer3_out_1130_U.if_read & AESL_inst_myproject.layer3_out_1130_U.if_empty_n;
    assign fifo_intf_2483.wr_en = AESL_inst_myproject.layer3_out_1130_U.if_write & AESL_inst_myproject.layer3_out_1130_U.if_full_n;
    assign fifo_intf_2483.fifo_rd_block = 0;
    assign fifo_intf_2483.fifo_wr_block = 0;
    assign fifo_intf_2483.finish = finish;
    csv_file_dump fifo_csv_dumper_2483;
    csv_file_dump cstatus_csv_dumper_2483;
    df_fifo_monitor fifo_monitor_2483;
    df_fifo_intf fifo_intf_2484(clock,reset);
    assign fifo_intf_2484.rd_en = AESL_inst_myproject.layer3_out_1131_U.if_read & AESL_inst_myproject.layer3_out_1131_U.if_empty_n;
    assign fifo_intf_2484.wr_en = AESL_inst_myproject.layer3_out_1131_U.if_write & AESL_inst_myproject.layer3_out_1131_U.if_full_n;
    assign fifo_intf_2484.fifo_rd_block = 0;
    assign fifo_intf_2484.fifo_wr_block = 0;
    assign fifo_intf_2484.finish = finish;
    csv_file_dump fifo_csv_dumper_2484;
    csv_file_dump cstatus_csv_dumper_2484;
    df_fifo_monitor fifo_monitor_2484;
    df_fifo_intf fifo_intf_2485(clock,reset);
    assign fifo_intf_2485.rd_en = AESL_inst_myproject.layer3_out_1132_U.if_read & AESL_inst_myproject.layer3_out_1132_U.if_empty_n;
    assign fifo_intf_2485.wr_en = AESL_inst_myproject.layer3_out_1132_U.if_write & AESL_inst_myproject.layer3_out_1132_U.if_full_n;
    assign fifo_intf_2485.fifo_rd_block = 0;
    assign fifo_intf_2485.fifo_wr_block = 0;
    assign fifo_intf_2485.finish = finish;
    csv_file_dump fifo_csv_dumper_2485;
    csv_file_dump cstatus_csv_dumper_2485;
    df_fifo_monitor fifo_monitor_2485;
    df_fifo_intf fifo_intf_2486(clock,reset);
    assign fifo_intf_2486.rd_en = AESL_inst_myproject.layer3_out_1133_U.if_read & AESL_inst_myproject.layer3_out_1133_U.if_empty_n;
    assign fifo_intf_2486.wr_en = AESL_inst_myproject.layer3_out_1133_U.if_write & AESL_inst_myproject.layer3_out_1133_U.if_full_n;
    assign fifo_intf_2486.fifo_rd_block = 0;
    assign fifo_intf_2486.fifo_wr_block = 0;
    assign fifo_intf_2486.finish = finish;
    csv_file_dump fifo_csv_dumper_2486;
    csv_file_dump cstatus_csv_dumper_2486;
    df_fifo_monitor fifo_monitor_2486;
    df_fifo_intf fifo_intf_2487(clock,reset);
    assign fifo_intf_2487.rd_en = AESL_inst_myproject.layer3_out_1134_U.if_read & AESL_inst_myproject.layer3_out_1134_U.if_empty_n;
    assign fifo_intf_2487.wr_en = AESL_inst_myproject.layer3_out_1134_U.if_write & AESL_inst_myproject.layer3_out_1134_U.if_full_n;
    assign fifo_intf_2487.fifo_rd_block = 0;
    assign fifo_intf_2487.fifo_wr_block = 0;
    assign fifo_intf_2487.finish = finish;
    csv_file_dump fifo_csv_dumper_2487;
    csv_file_dump cstatus_csv_dumper_2487;
    df_fifo_monitor fifo_monitor_2487;
    df_fifo_intf fifo_intf_2488(clock,reset);
    assign fifo_intf_2488.rd_en = AESL_inst_myproject.layer3_out_1135_U.if_read & AESL_inst_myproject.layer3_out_1135_U.if_empty_n;
    assign fifo_intf_2488.wr_en = AESL_inst_myproject.layer3_out_1135_U.if_write & AESL_inst_myproject.layer3_out_1135_U.if_full_n;
    assign fifo_intf_2488.fifo_rd_block = 0;
    assign fifo_intf_2488.fifo_wr_block = 0;
    assign fifo_intf_2488.finish = finish;
    csv_file_dump fifo_csv_dumper_2488;
    csv_file_dump cstatus_csv_dumper_2488;
    df_fifo_monitor fifo_monitor_2488;
    df_fifo_intf fifo_intf_2489(clock,reset);
    assign fifo_intf_2489.rd_en = AESL_inst_myproject.layer3_out_1136_U.if_read & AESL_inst_myproject.layer3_out_1136_U.if_empty_n;
    assign fifo_intf_2489.wr_en = AESL_inst_myproject.layer3_out_1136_U.if_write & AESL_inst_myproject.layer3_out_1136_U.if_full_n;
    assign fifo_intf_2489.fifo_rd_block = 0;
    assign fifo_intf_2489.fifo_wr_block = 0;
    assign fifo_intf_2489.finish = finish;
    csv_file_dump fifo_csv_dumper_2489;
    csv_file_dump cstatus_csv_dumper_2489;
    df_fifo_monitor fifo_monitor_2489;
    df_fifo_intf fifo_intf_2490(clock,reset);
    assign fifo_intf_2490.rd_en = AESL_inst_myproject.layer3_out_1137_U.if_read & AESL_inst_myproject.layer3_out_1137_U.if_empty_n;
    assign fifo_intf_2490.wr_en = AESL_inst_myproject.layer3_out_1137_U.if_write & AESL_inst_myproject.layer3_out_1137_U.if_full_n;
    assign fifo_intf_2490.fifo_rd_block = 0;
    assign fifo_intf_2490.fifo_wr_block = 0;
    assign fifo_intf_2490.finish = finish;
    csv_file_dump fifo_csv_dumper_2490;
    csv_file_dump cstatus_csv_dumper_2490;
    df_fifo_monitor fifo_monitor_2490;
    df_fifo_intf fifo_intf_2491(clock,reset);
    assign fifo_intf_2491.rd_en = AESL_inst_myproject.layer3_out_1138_U.if_read & AESL_inst_myproject.layer3_out_1138_U.if_empty_n;
    assign fifo_intf_2491.wr_en = AESL_inst_myproject.layer3_out_1138_U.if_write & AESL_inst_myproject.layer3_out_1138_U.if_full_n;
    assign fifo_intf_2491.fifo_rd_block = 0;
    assign fifo_intf_2491.fifo_wr_block = 0;
    assign fifo_intf_2491.finish = finish;
    csv_file_dump fifo_csv_dumper_2491;
    csv_file_dump cstatus_csv_dumper_2491;
    df_fifo_monitor fifo_monitor_2491;
    df_fifo_intf fifo_intf_2492(clock,reset);
    assign fifo_intf_2492.rd_en = AESL_inst_myproject.layer3_out_1139_U.if_read & AESL_inst_myproject.layer3_out_1139_U.if_empty_n;
    assign fifo_intf_2492.wr_en = AESL_inst_myproject.layer3_out_1139_U.if_write & AESL_inst_myproject.layer3_out_1139_U.if_full_n;
    assign fifo_intf_2492.fifo_rd_block = 0;
    assign fifo_intf_2492.fifo_wr_block = 0;
    assign fifo_intf_2492.finish = finish;
    csv_file_dump fifo_csv_dumper_2492;
    csv_file_dump cstatus_csv_dumper_2492;
    df_fifo_monitor fifo_monitor_2492;
    df_fifo_intf fifo_intf_2493(clock,reset);
    assign fifo_intf_2493.rd_en = AESL_inst_myproject.layer3_out_1140_U.if_read & AESL_inst_myproject.layer3_out_1140_U.if_empty_n;
    assign fifo_intf_2493.wr_en = AESL_inst_myproject.layer3_out_1140_U.if_write & AESL_inst_myproject.layer3_out_1140_U.if_full_n;
    assign fifo_intf_2493.fifo_rd_block = 0;
    assign fifo_intf_2493.fifo_wr_block = 0;
    assign fifo_intf_2493.finish = finish;
    csv_file_dump fifo_csv_dumper_2493;
    csv_file_dump cstatus_csv_dumper_2493;
    df_fifo_monitor fifo_monitor_2493;
    df_fifo_intf fifo_intf_2494(clock,reset);
    assign fifo_intf_2494.rd_en = AESL_inst_myproject.layer3_out_1141_U.if_read & AESL_inst_myproject.layer3_out_1141_U.if_empty_n;
    assign fifo_intf_2494.wr_en = AESL_inst_myproject.layer3_out_1141_U.if_write & AESL_inst_myproject.layer3_out_1141_U.if_full_n;
    assign fifo_intf_2494.fifo_rd_block = 0;
    assign fifo_intf_2494.fifo_wr_block = 0;
    assign fifo_intf_2494.finish = finish;
    csv_file_dump fifo_csv_dumper_2494;
    csv_file_dump cstatus_csv_dumper_2494;
    df_fifo_monitor fifo_monitor_2494;
    df_fifo_intf fifo_intf_2495(clock,reset);
    assign fifo_intf_2495.rd_en = AESL_inst_myproject.layer3_out_1142_U.if_read & AESL_inst_myproject.layer3_out_1142_U.if_empty_n;
    assign fifo_intf_2495.wr_en = AESL_inst_myproject.layer3_out_1142_U.if_write & AESL_inst_myproject.layer3_out_1142_U.if_full_n;
    assign fifo_intf_2495.fifo_rd_block = 0;
    assign fifo_intf_2495.fifo_wr_block = 0;
    assign fifo_intf_2495.finish = finish;
    csv_file_dump fifo_csv_dumper_2495;
    csv_file_dump cstatus_csv_dumper_2495;
    df_fifo_monitor fifo_monitor_2495;
    df_fifo_intf fifo_intf_2496(clock,reset);
    assign fifo_intf_2496.rd_en = AESL_inst_myproject.layer3_out_1143_U.if_read & AESL_inst_myproject.layer3_out_1143_U.if_empty_n;
    assign fifo_intf_2496.wr_en = AESL_inst_myproject.layer3_out_1143_U.if_write & AESL_inst_myproject.layer3_out_1143_U.if_full_n;
    assign fifo_intf_2496.fifo_rd_block = 0;
    assign fifo_intf_2496.fifo_wr_block = 0;
    assign fifo_intf_2496.finish = finish;
    csv_file_dump fifo_csv_dumper_2496;
    csv_file_dump cstatus_csv_dumper_2496;
    df_fifo_monitor fifo_monitor_2496;
    df_fifo_intf fifo_intf_2497(clock,reset);
    assign fifo_intf_2497.rd_en = AESL_inst_myproject.layer3_out_1144_U.if_read & AESL_inst_myproject.layer3_out_1144_U.if_empty_n;
    assign fifo_intf_2497.wr_en = AESL_inst_myproject.layer3_out_1144_U.if_write & AESL_inst_myproject.layer3_out_1144_U.if_full_n;
    assign fifo_intf_2497.fifo_rd_block = 0;
    assign fifo_intf_2497.fifo_wr_block = 0;
    assign fifo_intf_2497.finish = finish;
    csv_file_dump fifo_csv_dumper_2497;
    csv_file_dump cstatus_csv_dumper_2497;
    df_fifo_monitor fifo_monitor_2497;
    df_fifo_intf fifo_intf_2498(clock,reset);
    assign fifo_intf_2498.rd_en = AESL_inst_myproject.layer3_out_1145_U.if_read & AESL_inst_myproject.layer3_out_1145_U.if_empty_n;
    assign fifo_intf_2498.wr_en = AESL_inst_myproject.layer3_out_1145_U.if_write & AESL_inst_myproject.layer3_out_1145_U.if_full_n;
    assign fifo_intf_2498.fifo_rd_block = 0;
    assign fifo_intf_2498.fifo_wr_block = 0;
    assign fifo_intf_2498.finish = finish;
    csv_file_dump fifo_csv_dumper_2498;
    csv_file_dump cstatus_csv_dumper_2498;
    df_fifo_monitor fifo_monitor_2498;
    df_fifo_intf fifo_intf_2499(clock,reset);
    assign fifo_intf_2499.rd_en = AESL_inst_myproject.layer3_out_1146_U.if_read & AESL_inst_myproject.layer3_out_1146_U.if_empty_n;
    assign fifo_intf_2499.wr_en = AESL_inst_myproject.layer3_out_1146_U.if_write & AESL_inst_myproject.layer3_out_1146_U.if_full_n;
    assign fifo_intf_2499.fifo_rd_block = 0;
    assign fifo_intf_2499.fifo_wr_block = 0;
    assign fifo_intf_2499.finish = finish;
    csv_file_dump fifo_csv_dumper_2499;
    csv_file_dump cstatus_csv_dumper_2499;
    df_fifo_monitor fifo_monitor_2499;
    df_fifo_intf fifo_intf_2500(clock,reset);
    assign fifo_intf_2500.rd_en = AESL_inst_myproject.layer3_out_1147_U.if_read & AESL_inst_myproject.layer3_out_1147_U.if_empty_n;
    assign fifo_intf_2500.wr_en = AESL_inst_myproject.layer3_out_1147_U.if_write & AESL_inst_myproject.layer3_out_1147_U.if_full_n;
    assign fifo_intf_2500.fifo_rd_block = 0;
    assign fifo_intf_2500.fifo_wr_block = 0;
    assign fifo_intf_2500.finish = finish;
    csv_file_dump fifo_csv_dumper_2500;
    csv_file_dump cstatus_csv_dumper_2500;
    df_fifo_monitor fifo_monitor_2500;
    df_fifo_intf fifo_intf_2501(clock,reset);
    assign fifo_intf_2501.rd_en = AESL_inst_myproject.layer3_out_1148_U.if_read & AESL_inst_myproject.layer3_out_1148_U.if_empty_n;
    assign fifo_intf_2501.wr_en = AESL_inst_myproject.layer3_out_1148_U.if_write & AESL_inst_myproject.layer3_out_1148_U.if_full_n;
    assign fifo_intf_2501.fifo_rd_block = 0;
    assign fifo_intf_2501.fifo_wr_block = 0;
    assign fifo_intf_2501.finish = finish;
    csv_file_dump fifo_csv_dumper_2501;
    csv_file_dump cstatus_csv_dumper_2501;
    df_fifo_monitor fifo_monitor_2501;
    df_fifo_intf fifo_intf_2502(clock,reset);
    assign fifo_intf_2502.rd_en = AESL_inst_myproject.layer3_out_1149_U.if_read & AESL_inst_myproject.layer3_out_1149_U.if_empty_n;
    assign fifo_intf_2502.wr_en = AESL_inst_myproject.layer3_out_1149_U.if_write & AESL_inst_myproject.layer3_out_1149_U.if_full_n;
    assign fifo_intf_2502.fifo_rd_block = 0;
    assign fifo_intf_2502.fifo_wr_block = 0;
    assign fifo_intf_2502.finish = finish;
    csv_file_dump fifo_csv_dumper_2502;
    csv_file_dump cstatus_csv_dumper_2502;
    df_fifo_monitor fifo_monitor_2502;
    df_fifo_intf fifo_intf_2503(clock,reset);
    assign fifo_intf_2503.rd_en = AESL_inst_myproject.layer3_out_1150_U.if_read & AESL_inst_myproject.layer3_out_1150_U.if_empty_n;
    assign fifo_intf_2503.wr_en = AESL_inst_myproject.layer3_out_1150_U.if_write & AESL_inst_myproject.layer3_out_1150_U.if_full_n;
    assign fifo_intf_2503.fifo_rd_block = 0;
    assign fifo_intf_2503.fifo_wr_block = 0;
    assign fifo_intf_2503.finish = finish;
    csv_file_dump fifo_csv_dumper_2503;
    csv_file_dump cstatus_csv_dumper_2503;
    df_fifo_monitor fifo_monitor_2503;
    df_fifo_intf fifo_intf_2504(clock,reset);
    assign fifo_intf_2504.rd_en = AESL_inst_myproject.layer3_out_1151_U.if_read & AESL_inst_myproject.layer3_out_1151_U.if_empty_n;
    assign fifo_intf_2504.wr_en = AESL_inst_myproject.layer3_out_1151_U.if_write & AESL_inst_myproject.layer3_out_1151_U.if_full_n;
    assign fifo_intf_2504.fifo_rd_block = 0;
    assign fifo_intf_2504.fifo_wr_block = 0;
    assign fifo_intf_2504.finish = finish;
    csv_file_dump fifo_csv_dumper_2504;
    csv_file_dump cstatus_csv_dumper_2504;
    df_fifo_monitor fifo_monitor_2504;
    df_fifo_intf fifo_intf_2505(clock,reset);
    assign fifo_intf_2505.rd_en = AESL_inst_myproject.layer3_out_1152_U.if_read & AESL_inst_myproject.layer3_out_1152_U.if_empty_n;
    assign fifo_intf_2505.wr_en = AESL_inst_myproject.layer3_out_1152_U.if_write & AESL_inst_myproject.layer3_out_1152_U.if_full_n;
    assign fifo_intf_2505.fifo_rd_block = 0;
    assign fifo_intf_2505.fifo_wr_block = 0;
    assign fifo_intf_2505.finish = finish;
    csv_file_dump fifo_csv_dumper_2505;
    csv_file_dump cstatus_csv_dumper_2505;
    df_fifo_monitor fifo_monitor_2505;
    df_fifo_intf fifo_intf_2506(clock,reset);
    assign fifo_intf_2506.rd_en = AESL_inst_myproject.layer3_out_1153_U.if_read & AESL_inst_myproject.layer3_out_1153_U.if_empty_n;
    assign fifo_intf_2506.wr_en = AESL_inst_myproject.layer3_out_1153_U.if_write & AESL_inst_myproject.layer3_out_1153_U.if_full_n;
    assign fifo_intf_2506.fifo_rd_block = 0;
    assign fifo_intf_2506.fifo_wr_block = 0;
    assign fifo_intf_2506.finish = finish;
    csv_file_dump fifo_csv_dumper_2506;
    csv_file_dump cstatus_csv_dumper_2506;
    df_fifo_monitor fifo_monitor_2506;
    df_fifo_intf fifo_intf_2507(clock,reset);
    assign fifo_intf_2507.rd_en = AESL_inst_myproject.layer3_out_1154_U.if_read & AESL_inst_myproject.layer3_out_1154_U.if_empty_n;
    assign fifo_intf_2507.wr_en = AESL_inst_myproject.layer3_out_1154_U.if_write & AESL_inst_myproject.layer3_out_1154_U.if_full_n;
    assign fifo_intf_2507.fifo_rd_block = 0;
    assign fifo_intf_2507.fifo_wr_block = 0;
    assign fifo_intf_2507.finish = finish;
    csv_file_dump fifo_csv_dumper_2507;
    csv_file_dump cstatus_csv_dumper_2507;
    df_fifo_monitor fifo_monitor_2507;
    df_fifo_intf fifo_intf_2508(clock,reset);
    assign fifo_intf_2508.rd_en = AESL_inst_myproject.layer3_out_1155_U.if_read & AESL_inst_myproject.layer3_out_1155_U.if_empty_n;
    assign fifo_intf_2508.wr_en = AESL_inst_myproject.layer3_out_1155_U.if_write & AESL_inst_myproject.layer3_out_1155_U.if_full_n;
    assign fifo_intf_2508.fifo_rd_block = 0;
    assign fifo_intf_2508.fifo_wr_block = 0;
    assign fifo_intf_2508.finish = finish;
    csv_file_dump fifo_csv_dumper_2508;
    csv_file_dump cstatus_csv_dumper_2508;
    df_fifo_monitor fifo_monitor_2508;
    df_fifo_intf fifo_intf_2509(clock,reset);
    assign fifo_intf_2509.rd_en = AESL_inst_myproject.layer3_out_1156_U.if_read & AESL_inst_myproject.layer3_out_1156_U.if_empty_n;
    assign fifo_intf_2509.wr_en = AESL_inst_myproject.layer3_out_1156_U.if_write & AESL_inst_myproject.layer3_out_1156_U.if_full_n;
    assign fifo_intf_2509.fifo_rd_block = 0;
    assign fifo_intf_2509.fifo_wr_block = 0;
    assign fifo_intf_2509.finish = finish;
    csv_file_dump fifo_csv_dumper_2509;
    csv_file_dump cstatus_csv_dumper_2509;
    df_fifo_monitor fifo_monitor_2509;
    df_fifo_intf fifo_intf_2510(clock,reset);
    assign fifo_intf_2510.rd_en = AESL_inst_myproject.layer3_out_1157_U.if_read & AESL_inst_myproject.layer3_out_1157_U.if_empty_n;
    assign fifo_intf_2510.wr_en = AESL_inst_myproject.layer3_out_1157_U.if_write & AESL_inst_myproject.layer3_out_1157_U.if_full_n;
    assign fifo_intf_2510.fifo_rd_block = 0;
    assign fifo_intf_2510.fifo_wr_block = 0;
    assign fifo_intf_2510.finish = finish;
    csv_file_dump fifo_csv_dumper_2510;
    csv_file_dump cstatus_csv_dumper_2510;
    df_fifo_monitor fifo_monitor_2510;
    df_fifo_intf fifo_intf_2511(clock,reset);
    assign fifo_intf_2511.rd_en = AESL_inst_myproject.layer3_out_1158_U.if_read & AESL_inst_myproject.layer3_out_1158_U.if_empty_n;
    assign fifo_intf_2511.wr_en = AESL_inst_myproject.layer3_out_1158_U.if_write & AESL_inst_myproject.layer3_out_1158_U.if_full_n;
    assign fifo_intf_2511.fifo_rd_block = 0;
    assign fifo_intf_2511.fifo_wr_block = 0;
    assign fifo_intf_2511.finish = finish;
    csv_file_dump fifo_csv_dumper_2511;
    csv_file_dump cstatus_csv_dumper_2511;
    df_fifo_monitor fifo_monitor_2511;
    df_fifo_intf fifo_intf_2512(clock,reset);
    assign fifo_intf_2512.rd_en = AESL_inst_myproject.layer3_out_1159_U.if_read & AESL_inst_myproject.layer3_out_1159_U.if_empty_n;
    assign fifo_intf_2512.wr_en = AESL_inst_myproject.layer3_out_1159_U.if_write & AESL_inst_myproject.layer3_out_1159_U.if_full_n;
    assign fifo_intf_2512.fifo_rd_block = 0;
    assign fifo_intf_2512.fifo_wr_block = 0;
    assign fifo_intf_2512.finish = finish;
    csv_file_dump fifo_csv_dumper_2512;
    csv_file_dump cstatus_csv_dumper_2512;
    df_fifo_monitor fifo_monitor_2512;
    df_fifo_intf fifo_intf_2513(clock,reset);
    assign fifo_intf_2513.rd_en = AESL_inst_myproject.layer3_out_1160_U.if_read & AESL_inst_myproject.layer3_out_1160_U.if_empty_n;
    assign fifo_intf_2513.wr_en = AESL_inst_myproject.layer3_out_1160_U.if_write & AESL_inst_myproject.layer3_out_1160_U.if_full_n;
    assign fifo_intf_2513.fifo_rd_block = 0;
    assign fifo_intf_2513.fifo_wr_block = 0;
    assign fifo_intf_2513.finish = finish;
    csv_file_dump fifo_csv_dumper_2513;
    csv_file_dump cstatus_csv_dumper_2513;
    df_fifo_monitor fifo_monitor_2513;
    df_fifo_intf fifo_intf_2514(clock,reset);
    assign fifo_intf_2514.rd_en = AESL_inst_myproject.layer3_out_1161_U.if_read & AESL_inst_myproject.layer3_out_1161_U.if_empty_n;
    assign fifo_intf_2514.wr_en = AESL_inst_myproject.layer3_out_1161_U.if_write & AESL_inst_myproject.layer3_out_1161_U.if_full_n;
    assign fifo_intf_2514.fifo_rd_block = 0;
    assign fifo_intf_2514.fifo_wr_block = 0;
    assign fifo_intf_2514.finish = finish;
    csv_file_dump fifo_csv_dumper_2514;
    csv_file_dump cstatus_csv_dumper_2514;
    df_fifo_monitor fifo_monitor_2514;
    df_fifo_intf fifo_intf_2515(clock,reset);
    assign fifo_intf_2515.rd_en = AESL_inst_myproject.layer3_out_1162_U.if_read & AESL_inst_myproject.layer3_out_1162_U.if_empty_n;
    assign fifo_intf_2515.wr_en = AESL_inst_myproject.layer3_out_1162_U.if_write & AESL_inst_myproject.layer3_out_1162_U.if_full_n;
    assign fifo_intf_2515.fifo_rd_block = 0;
    assign fifo_intf_2515.fifo_wr_block = 0;
    assign fifo_intf_2515.finish = finish;
    csv_file_dump fifo_csv_dumper_2515;
    csv_file_dump cstatus_csv_dumper_2515;
    df_fifo_monitor fifo_monitor_2515;
    df_fifo_intf fifo_intf_2516(clock,reset);
    assign fifo_intf_2516.rd_en = AESL_inst_myproject.layer3_out_1163_U.if_read & AESL_inst_myproject.layer3_out_1163_U.if_empty_n;
    assign fifo_intf_2516.wr_en = AESL_inst_myproject.layer3_out_1163_U.if_write & AESL_inst_myproject.layer3_out_1163_U.if_full_n;
    assign fifo_intf_2516.fifo_rd_block = 0;
    assign fifo_intf_2516.fifo_wr_block = 0;
    assign fifo_intf_2516.finish = finish;
    csv_file_dump fifo_csv_dumper_2516;
    csv_file_dump cstatus_csv_dumper_2516;
    df_fifo_monitor fifo_monitor_2516;
    df_fifo_intf fifo_intf_2517(clock,reset);
    assign fifo_intf_2517.rd_en = AESL_inst_myproject.layer3_out_1164_U.if_read & AESL_inst_myproject.layer3_out_1164_U.if_empty_n;
    assign fifo_intf_2517.wr_en = AESL_inst_myproject.layer3_out_1164_U.if_write & AESL_inst_myproject.layer3_out_1164_U.if_full_n;
    assign fifo_intf_2517.fifo_rd_block = 0;
    assign fifo_intf_2517.fifo_wr_block = 0;
    assign fifo_intf_2517.finish = finish;
    csv_file_dump fifo_csv_dumper_2517;
    csv_file_dump cstatus_csv_dumper_2517;
    df_fifo_monitor fifo_monitor_2517;
    df_fifo_intf fifo_intf_2518(clock,reset);
    assign fifo_intf_2518.rd_en = AESL_inst_myproject.layer3_out_1165_U.if_read & AESL_inst_myproject.layer3_out_1165_U.if_empty_n;
    assign fifo_intf_2518.wr_en = AESL_inst_myproject.layer3_out_1165_U.if_write & AESL_inst_myproject.layer3_out_1165_U.if_full_n;
    assign fifo_intf_2518.fifo_rd_block = 0;
    assign fifo_intf_2518.fifo_wr_block = 0;
    assign fifo_intf_2518.finish = finish;
    csv_file_dump fifo_csv_dumper_2518;
    csv_file_dump cstatus_csv_dumper_2518;
    df_fifo_monitor fifo_monitor_2518;
    df_fifo_intf fifo_intf_2519(clock,reset);
    assign fifo_intf_2519.rd_en = AESL_inst_myproject.layer3_out_1166_U.if_read & AESL_inst_myproject.layer3_out_1166_U.if_empty_n;
    assign fifo_intf_2519.wr_en = AESL_inst_myproject.layer3_out_1166_U.if_write & AESL_inst_myproject.layer3_out_1166_U.if_full_n;
    assign fifo_intf_2519.fifo_rd_block = 0;
    assign fifo_intf_2519.fifo_wr_block = 0;
    assign fifo_intf_2519.finish = finish;
    csv_file_dump fifo_csv_dumper_2519;
    csv_file_dump cstatus_csv_dumper_2519;
    df_fifo_monitor fifo_monitor_2519;
    df_fifo_intf fifo_intf_2520(clock,reset);
    assign fifo_intf_2520.rd_en = AESL_inst_myproject.layer3_out_1167_U.if_read & AESL_inst_myproject.layer3_out_1167_U.if_empty_n;
    assign fifo_intf_2520.wr_en = AESL_inst_myproject.layer3_out_1167_U.if_write & AESL_inst_myproject.layer3_out_1167_U.if_full_n;
    assign fifo_intf_2520.fifo_rd_block = 0;
    assign fifo_intf_2520.fifo_wr_block = 0;
    assign fifo_intf_2520.finish = finish;
    csv_file_dump fifo_csv_dumper_2520;
    csv_file_dump cstatus_csv_dumper_2520;
    df_fifo_monitor fifo_monitor_2520;
    df_fifo_intf fifo_intf_2521(clock,reset);
    assign fifo_intf_2521.rd_en = AESL_inst_myproject.layer3_out_1168_U.if_read & AESL_inst_myproject.layer3_out_1168_U.if_empty_n;
    assign fifo_intf_2521.wr_en = AESL_inst_myproject.layer3_out_1168_U.if_write & AESL_inst_myproject.layer3_out_1168_U.if_full_n;
    assign fifo_intf_2521.fifo_rd_block = 0;
    assign fifo_intf_2521.fifo_wr_block = 0;
    assign fifo_intf_2521.finish = finish;
    csv_file_dump fifo_csv_dumper_2521;
    csv_file_dump cstatus_csv_dumper_2521;
    df_fifo_monitor fifo_monitor_2521;
    df_fifo_intf fifo_intf_2522(clock,reset);
    assign fifo_intf_2522.rd_en = AESL_inst_myproject.layer3_out_1169_U.if_read & AESL_inst_myproject.layer3_out_1169_U.if_empty_n;
    assign fifo_intf_2522.wr_en = AESL_inst_myproject.layer3_out_1169_U.if_write & AESL_inst_myproject.layer3_out_1169_U.if_full_n;
    assign fifo_intf_2522.fifo_rd_block = 0;
    assign fifo_intf_2522.fifo_wr_block = 0;
    assign fifo_intf_2522.finish = finish;
    csv_file_dump fifo_csv_dumper_2522;
    csv_file_dump cstatus_csv_dumper_2522;
    df_fifo_monitor fifo_monitor_2522;
    df_fifo_intf fifo_intf_2523(clock,reset);
    assign fifo_intf_2523.rd_en = AESL_inst_myproject.layer3_out_1170_U.if_read & AESL_inst_myproject.layer3_out_1170_U.if_empty_n;
    assign fifo_intf_2523.wr_en = AESL_inst_myproject.layer3_out_1170_U.if_write & AESL_inst_myproject.layer3_out_1170_U.if_full_n;
    assign fifo_intf_2523.fifo_rd_block = 0;
    assign fifo_intf_2523.fifo_wr_block = 0;
    assign fifo_intf_2523.finish = finish;
    csv_file_dump fifo_csv_dumper_2523;
    csv_file_dump cstatus_csv_dumper_2523;
    df_fifo_monitor fifo_monitor_2523;
    df_fifo_intf fifo_intf_2524(clock,reset);
    assign fifo_intf_2524.rd_en = AESL_inst_myproject.layer3_out_1171_U.if_read & AESL_inst_myproject.layer3_out_1171_U.if_empty_n;
    assign fifo_intf_2524.wr_en = AESL_inst_myproject.layer3_out_1171_U.if_write & AESL_inst_myproject.layer3_out_1171_U.if_full_n;
    assign fifo_intf_2524.fifo_rd_block = 0;
    assign fifo_intf_2524.fifo_wr_block = 0;
    assign fifo_intf_2524.finish = finish;
    csv_file_dump fifo_csv_dumper_2524;
    csv_file_dump cstatus_csv_dumper_2524;
    df_fifo_monitor fifo_monitor_2524;
    df_fifo_intf fifo_intf_2525(clock,reset);
    assign fifo_intf_2525.rd_en = AESL_inst_myproject.layer3_out_1172_U.if_read & AESL_inst_myproject.layer3_out_1172_U.if_empty_n;
    assign fifo_intf_2525.wr_en = AESL_inst_myproject.layer3_out_1172_U.if_write & AESL_inst_myproject.layer3_out_1172_U.if_full_n;
    assign fifo_intf_2525.fifo_rd_block = 0;
    assign fifo_intf_2525.fifo_wr_block = 0;
    assign fifo_intf_2525.finish = finish;
    csv_file_dump fifo_csv_dumper_2525;
    csv_file_dump cstatus_csv_dumper_2525;
    df_fifo_monitor fifo_monitor_2525;
    df_fifo_intf fifo_intf_2526(clock,reset);
    assign fifo_intf_2526.rd_en = AESL_inst_myproject.layer3_out_1173_U.if_read & AESL_inst_myproject.layer3_out_1173_U.if_empty_n;
    assign fifo_intf_2526.wr_en = AESL_inst_myproject.layer3_out_1173_U.if_write & AESL_inst_myproject.layer3_out_1173_U.if_full_n;
    assign fifo_intf_2526.fifo_rd_block = 0;
    assign fifo_intf_2526.fifo_wr_block = 0;
    assign fifo_intf_2526.finish = finish;
    csv_file_dump fifo_csv_dumper_2526;
    csv_file_dump cstatus_csv_dumper_2526;
    df_fifo_monitor fifo_monitor_2526;
    df_fifo_intf fifo_intf_2527(clock,reset);
    assign fifo_intf_2527.rd_en = AESL_inst_myproject.layer3_out_1174_U.if_read & AESL_inst_myproject.layer3_out_1174_U.if_empty_n;
    assign fifo_intf_2527.wr_en = AESL_inst_myproject.layer3_out_1174_U.if_write & AESL_inst_myproject.layer3_out_1174_U.if_full_n;
    assign fifo_intf_2527.fifo_rd_block = 0;
    assign fifo_intf_2527.fifo_wr_block = 0;
    assign fifo_intf_2527.finish = finish;
    csv_file_dump fifo_csv_dumper_2527;
    csv_file_dump cstatus_csv_dumper_2527;
    df_fifo_monitor fifo_monitor_2527;
    df_fifo_intf fifo_intf_2528(clock,reset);
    assign fifo_intf_2528.rd_en = AESL_inst_myproject.layer3_out_1175_U.if_read & AESL_inst_myproject.layer3_out_1175_U.if_empty_n;
    assign fifo_intf_2528.wr_en = AESL_inst_myproject.layer3_out_1175_U.if_write & AESL_inst_myproject.layer3_out_1175_U.if_full_n;
    assign fifo_intf_2528.fifo_rd_block = 0;
    assign fifo_intf_2528.fifo_wr_block = 0;
    assign fifo_intf_2528.finish = finish;
    csv_file_dump fifo_csv_dumper_2528;
    csv_file_dump cstatus_csv_dumper_2528;
    df_fifo_monitor fifo_monitor_2528;
    df_fifo_intf fifo_intf_2529(clock,reset);
    assign fifo_intf_2529.rd_en = AESL_inst_myproject.layer3_out_1176_U.if_read & AESL_inst_myproject.layer3_out_1176_U.if_empty_n;
    assign fifo_intf_2529.wr_en = AESL_inst_myproject.layer3_out_1176_U.if_write & AESL_inst_myproject.layer3_out_1176_U.if_full_n;
    assign fifo_intf_2529.fifo_rd_block = 0;
    assign fifo_intf_2529.fifo_wr_block = 0;
    assign fifo_intf_2529.finish = finish;
    csv_file_dump fifo_csv_dumper_2529;
    csv_file_dump cstatus_csv_dumper_2529;
    df_fifo_monitor fifo_monitor_2529;
    df_fifo_intf fifo_intf_2530(clock,reset);
    assign fifo_intf_2530.rd_en = AESL_inst_myproject.layer3_out_1177_U.if_read & AESL_inst_myproject.layer3_out_1177_U.if_empty_n;
    assign fifo_intf_2530.wr_en = AESL_inst_myproject.layer3_out_1177_U.if_write & AESL_inst_myproject.layer3_out_1177_U.if_full_n;
    assign fifo_intf_2530.fifo_rd_block = 0;
    assign fifo_intf_2530.fifo_wr_block = 0;
    assign fifo_intf_2530.finish = finish;
    csv_file_dump fifo_csv_dumper_2530;
    csv_file_dump cstatus_csv_dumper_2530;
    df_fifo_monitor fifo_monitor_2530;
    df_fifo_intf fifo_intf_2531(clock,reset);
    assign fifo_intf_2531.rd_en = AESL_inst_myproject.layer3_out_1178_U.if_read & AESL_inst_myproject.layer3_out_1178_U.if_empty_n;
    assign fifo_intf_2531.wr_en = AESL_inst_myproject.layer3_out_1178_U.if_write & AESL_inst_myproject.layer3_out_1178_U.if_full_n;
    assign fifo_intf_2531.fifo_rd_block = 0;
    assign fifo_intf_2531.fifo_wr_block = 0;
    assign fifo_intf_2531.finish = finish;
    csv_file_dump fifo_csv_dumper_2531;
    csv_file_dump cstatus_csv_dumper_2531;
    df_fifo_monitor fifo_monitor_2531;
    df_fifo_intf fifo_intf_2532(clock,reset);
    assign fifo_intf_2532.rd_en = AESL_inst_myproject.layer3_out_1179_U.if_read & AESL_inst_myproject.layer3_out_1179_U.if_empty_n;
    assign fifo_intf_2532.wr_en = AESL_inst_myproject.layer3_out_1179_U.if_write & AESL_inst_myproject.layer3_out_1179_U.if_full_n;
    assign fifo_intf_2532.fifo_rd_block = 0;
    assign fifo_intf_2532.fifo_wr_block = 0;
    assign fifo_intf_2532.finish = finish;
    csv_file_dump fifo_csv_dumper_2532;
    csv_file_dump cstatus_csv_dumper_2532;
    df_fifo_monitor fifo_monitor_2532;
    df_fifo_intf fifo_intf_2533(clock,reset);
    assign fifo_intf_2533.rd_en = AESL_inst_myproject.layer3_out_1180_U.if_read & AESL_inst_myproject.layer3_out_1180_U.if_empty_n;
    assign fifo_intf_2533.wr_en = AESL_inst_myproject.layer3_out_1180_U.if_write & AESL_inst_myproject.layer3_out_1180_U.if_full_n;
    assign fifo_intf_2533.fifo_rd_block = 0;
    assign fifo_intf_2533.fifo_wr_block = 0;
    assign fifo_intf_2533.finish = finish;
    csv_file_dump fifo_csv_dumper_2533;
    csv_file_dump cstatus_csv_dumper_2533;
    df_fifo_monitor fifo_monitor_2533;
    df_fifo_intf fifo_intf_2534(clock,reset);
    assign fifo_intf_2534.rd_en = AESL_inst_myproject.layer3_out_1181_U.if_read & AESL_inst_myproject.layer3_out_1181_U.if_empty_n;
    assign fifo_intf_2534.wr_en = AESL_inst_myproject.layer3_out_1181_U.if_write & AESL_inst_myproject.layer3_out_1181_U.if_full_n;
    assign fifo_intf_2534.fifo_rd_block = 0;
    assign fifo_intf_2534.fifo_wr_block = 0;
    assign fifo_intf_2534.finish = finish;
    csv_file_dump fifo_csv_dumper_2534;
    csv_file_dump cstatus_csv_dumper_2534;
    df_fifo_monitor fifo_monitor_2534;
    df_fifo_intf fifo_intf_2535(clock,reset);
    assign fifo_intf_2535.rd_en = AESL_inst_myproject.layer3_out_1182_U.if_read & AESL_inst_myproject.layer3_out_1182_U.if_empty_n;
    assign fifo_intf_2535.wr_en = AESL_inst_myproject.layer3_out_1182_U.if_write & AESL_inst_myproject.layer3_out_1182_U.if_full_n;
    assign fifo_intf_2535.fifo_rd_block = 0;
    assign fifo_intf_2535.fifo_wr_block = 0;
    assign fifo_intf_2535.finish = finish;
    csv_file_dump fifo_csv_dumper_2535;
    csv_file_dump cstatus_csv_dumper_2535;
    df_fifo_monitor fifo_monitor_2535;
    df_fifo_intf fifo_intf_2536(clock,reset);
    assign fifo_intf_2536.rd_en = AESL_inst_myproject.layer3_out_1183_U.if_read & AESL_inst_myproject.layer3_out_1183_U.if_empty_n;
    assign fifo_intf_2536.wr_en = AESL_inst_myproject.layer3_out_1183_U.if_write & AESL_inst_myproject.layer3_out_1183_U.if_full_n;
    assign fifo_intf_2536.fifo_rd_block = 0;
    assign fifo_intf_2536.fifo_wr_block = 0;
    assign fifo_intf_2536.finish = finish;
    csv_file_dump fifo_csv_dumper_2536;
    csv_file_dump cstatus_csv_dumper_2536;
    df_fifo_monitor fifo_monitor_2536;
    df_fifo_intf fifo_intf_2537(clock,reset);
    assign fifo_intf_2537.rd_en = AESL_inst_myproject.layer3_out_1184_U.if_read & AESL_inst_myproject.layer3_out_1184_U.if_empty_n;
    assign fifo_intf_2537.wr_en = AESL_inst_myproject.layer3_out_1184_U.if_write & AESL_inst_myproject.layer3_out_1184_U.if_full_n;
    assign fifo_intf_2537.fifo_rd_block = 0;
    assign fifo_intf_2537.fifo_wr_block = 0;
    assign fifo_intf_2537.finish = finish;
    csv_file_dump fifo_csv_dumper_2537;
    csv_file_dump cstatus_csv_dumper_2537;
    df_fifo_monitor fifo_monitor_2537;
    df_fifo_intf fifo_intf_2538(clock,reset);
    assign fifo_intf_2538.rd_en = AESL_inst_myproject.layer3_out_1185_U.if_read & AESL_inst_myproject.layer3_out_1185_U.if_empty_n;
    assign fifo_intf_2538.wr_en = AESL_inst_myproject.layer3_out_1185_U.if_write & AESL_inst_myproject.layer3_out_1185_U.if_full_n;
    assign fifo_intf_2538.fifo_rd_block = 0;
    assign fifo_intf_2538.fifo_wr_block = 0;
    assign fifo_intf_2538.finish = finish;
    csv_file_dump fifo_csv_dumper_2538;
    csv_file_dump cstatus_csv_dumper_2538;
    df_fifo_monitor fifo_monitor_2538;
    df_fifo_intf fifo_intf_2539(clock,reset);
    assign fifo_intf_2539.rd_en = AESL_inst_myproject.layer3_out_1186_U.if_read & AESL_inst_myproject.layer3_out_1186_U.if_empty_n;
    assign fifo_intf_2539.wr_en = AESL_inst_myproject.layer3_out_1186_U.if_write & AESL_inst_myproject.layer3_out_1186_U.if_full_n;
    assign fifo_intf_2539.fifo_rd_block = 0;
    assign fifo_intf_2539.fifo_wr_block = 0;
    assign fifo_intf_2539.finish = finish;
    csv_file_dump fifo_csv_dumper_2539;
    csv_file_dump cstatus_csv_dumper_2539;
    df_fifo_monitor fifo_monitor_2539;
    df_fifo_intf fifo_intf_2540(clock,reset);
    assign fifo_intf_2540.rd_en = AESL_inst_myproject.layer3_out_1187_U.if_read & AESL_inst_myproject.layer3_out_1187_U.if_empty_n;
    assign fifo_intf_2540.wr_en = AESL_inst_myproject.layer3_out_1187_U.if_write & AESL_inst_myproject.layer3_out_1187_U.if_full_n;
    assign fifo_intf_2540.fifo_rd_block = 0;
    assign fifo_intf_2540.fifo_wr_block = 0;
    assign fifo_intf_2540.finish = finish;
    csv_file_dump fifo_csv_dumper_2540;
    csv_file_dump cstatus_csv_dumper_2540;
    df_fifo_monitor fifo_monitor_2540;
    df_fifo_intf fifo_intf_2541(clock,reset);
    assign fifo_intf_2541.rd_en = AESL_inst_myproject.layer3_out_1188_U.if_read & AESL_inst_myproject.layer3_out_1188_U.if_empty_n;
    assign fifo_intf_2541.wr_en = AESL_inst_myproject.layer3_out_1188_U.if_write & AESL_inst_myproject.layer3_out_1188_U.if_full_n;
    assign fifo_intf_2541.fifo_rd_block = 0;
    assign fifo_intf_2541.fifo_wr_block = 0;
    assign fifo_intf_2541.finish = finish;
    csv_file_dump fifo_csv_dumper_2541;
    csv_file_dump cstatus_csv_dumper_2541;
    df_fifo_monitor fifo_monitor_2541;
    df_fifo_intf fifo_intf_2542(clock,reset);
    assign fifo_intf_2542.rd_en = AESL_inst_myproject.layer3_out_1189_U.if_read & AESL_inst_myproject.layer3_out_1189_U.if_empty_n;
    assign fifo_intf_2542.wr_en = AESL_inst_myproject.layer3_out_1189_U.if_write & AESL_inst_myproject.layer3_out_1189_U.if_full_n;
    assign fifo_intf_2542.fifo_rd_block = 0;
    assign fifo_intf_2542.fifo_wr_block = 0;
    assign fifo_intf_2542.finish = finish;
    csv_file_dump fifo_csv_dumper_2542;
    csv_file_dump cstatus_csv_dumper_2542;
    df_fifo_monitor fifo_monitor_2542;
    df_fifo_intf fifo_intf_2543(clock,reset);
    assign fifo_intf_2543.rd_en = AESL_inst_myproject.layer3_out_1190_U.if_read & AESL_inst_myproject.layer3_out_1190_U.if_empty_n;
    assign fifo_intf_2543.wr_en = AESL_inst_myproject.layer3_out_1190_U.if_write & AESL_inst_myproject.layer3_out_1190_U.if_full_n;
    assign fifo_intf_2543.fifo_rd_block = 0;
    assign fifo_intf_2543.fifo_wr_block = 0;
    assign fifo_intf_2543.finish = finish;
    csv_file_dump fifo_csv_dumper_2543;
    csv_file_dump cstatus_csv_dumper_2543;
    df_fifo_monitor fifo_monitor_2543;
    df_fifo_intf fifo_intf_2544(clock,reset);
    assign fifo_intf_2544.rd_en = AESL_inst_myproject.layer3_out_1191_U.if_read & AESL_inst_myproject.layer3_out_1191_U.if_empty_n;
    assign fifo_intf_2544.wr_en = AESL_inst_myproject.layer3_out_1191_U.if_write & AESL_inst_myproject.layer3_out_1191_U.if_full_n;
    assign fifo_intf_2544.fifo_rd_block = 0;
    assign fifo_intf_2544.fifo_wr_block = 0;
    assign fifo_intf_2544.finish = finish;
    csv_file_dump fifo_csv_dumper_2544;
    csv_file_dump cstatus_csv_dumper_2544;
    df_fifo_monitor fifo_monitor_2544;
    df_fifo_intf fifo_intf_2545(clock,reset);
    assign fifo_intf_2545.rd_en = AESL_inst_myproject.layer3_out_1192_U.if_read & AESL_inst_myproject.layer3_out_1192_U.if_empty_n;
    assign fifo_intf_2545.wr_en = AESL_inst_myproject.layer3_out_1192_U.if_write & AESL_inst_myproject.layer3_out_1192_U.if_full_n;
    assign fifo_intf_2545.fifo_rd_block = 0;
    assign fifo_intf_2545.fifo_wr_block = 0;
    assign fifo_intf_2545.finish = finish;
    csv_file_dump fifo_csv_dumper_2545;
    csv_file_dump cstatus_csv_dumper_2545;
    df_fifo_monitor fifo_monitor_2545;
    df_fifo_intf fifo_intf_2546(clock,reset);
    assign fifo_intf_2546.rd_en = AESL_inst_myproject.layer3_out_1193_U.if_read & AESL_inst_myproject.layer3_out_1193_U.if_empty_n;
    assign fifo_intf_2546.wr_en = AESL_inst_myproject.layer3_out_1193_U.if_write & AESL_inst_myproject.layer3_out_1193_U.if_full_n;
    assign fifo_intf_2546.fifo_rd_block = 0;
    assign fifo_intf_2546.fifo_wr_block = 0;
    assign fifo_intf_2546.finish = finish;
    csv_file_dump fifo_csv_dumper_2546;
    csv_file_dump cstatus_csv_dumper_2546;
    df_fifo_monitor fifo_monitor_2546;
    df_fifo_intf fifo_intf_2547(clock,reset);
    assign fifo_intf_2547.rd_en = AESL_inst_myproject.layer3_out_1194_U.if_read & AESL_inst_myproject.layer3_out_1194_U.if_empty_n;
    assign fifo_intf_2547.wr_en = AESL_inst_myproject.layer3_out_1194_U.if_write & AESL_inst_myproject.layer3_out_1194_U.if_full_n;
    assign fifo_intf_2547.fifo_rd_block = 0;
    assign fifo_intf_2547.fifo_wr_block = 0;
    assign fifo_intf_2547.finish = finish;
    csv_file_dump fifo_csv_dumper_2547;
    csv_file_dump cstatus_csv_dumper_2547;
    df_fifo_monitor fifo_monitor_2547;
    df_fifo_intf fifo_intf_2548(clock,reset);
    assign fifo_intf_2548.rd_en = AESL_inst_myproject.layer3_out_1195_U.if_read & AESL_inst_myproject.layer3_out_1195_U.if_empty_n;
    assign fifo_intf_2548.wr_en = AESL_inst_myproject.layer3_out_1195_U.if_write & AESL_inst_myproject.layer3_out_1195_U.if_full_n;
    assign fifo_intf_2548.fifo_rd_block = 0;
    assign fifo_intf_2548.fifo_wr_block = 0;
    assign fifo_intf_2548.finish = finish;
    csv_file_dump fifo_csv_dumper_2548;
    csv_file_dump cstatus_csv_dumper_2548;
    df_fifo_monitor fifo_monitor_2548;
    df_fifo_intf fifo_intf_2549(clock,reset);
    assign fifo_intf_2549.rd_en = AESL_inst_myproject.layer3_out_1196_U.if_read & AESL_inst_myproject.layer3_out_1196_U.if_empty_n;
    assign fifo_intf_2549.wr_en = AESL_inst_myproject.layer3_out_1196_U.if_write & AESL_inst_myproject.layer3_out_1196_U.if_full_n;
    assign fifo_intf_2549.fifo_rd_block = 0;
    assign fifo_intf_2549.fifo_wr_block = 0;
    assign fifo_intf_2549.finish = finish;
    csv_file_dump fifo_csv_dumper_2549;
    csv_file_dump cstatus_csv_dumper_2549;
    df_fifo_monitor fifo_monitor_2549;
    df_fifo_intf fifo_intf_2550(clock,reset);
    assign fifo_intf_2550.rd_en = AESL_inst_myproject.layer3_out_1197_U.if_read & AESL_inst_myproject.layer3_out_1197_U.if_empty_n;
    assign fifo_intf_2550.wr_en = AESL_inst_myproject.layer3_out_1197_U.if_write & AESL_inst_myproject.layer3_out_1197_U.if_full_n;
    assign fifo_intf_2550.fifo_rd_block = 0;
    assign fifo_intf_2550.fifo_wr_block = 0;
    assign fifo_intf_2550.finish = finish;
    csv_file_dump fifo_csv_dumper_2550;
    csv_file_dump cstatus_csv_dumper_2550;
    df_fifo_monitor fifo_monitor_2550;
    df_fifo_intf fifo_intf_2551(clock,reset);
    assign fifo_intf_2551.rd_en = AESL_inst_myproject.layer3_out_1198_U.if_read & AESL_inst_myproject.layer3_out_1198_U.if_empty_n;
    assign fifo_intf_2551.wr_en = AESL_inst_myproject.layer3_out_1198_U.if_write & AESL_inst_myproject.layer3_out_1198_U.if_full_n;
    assign fifo_intf_2551.fifo_rd_block = 0;
    assign fifo_intf_2551.fifo_wr_block = 0;
    assign fifo_intf_2551.finish = finish;
    csv_file_dump fifo_csv_dumper_2551;
    csv_file_dump cstatus_csv_dumper_2551;
    df_fifo_monitor fifo_monitor_2551;
    df_fifo_intf fifo_intf_2552(clock,reset);
    assign fifo_intf_2552.rd_en = AESL_inst_myproject.layer3_out_1199_U.if_read & AESL_inst_myproject.layer3_out_1199_U.if_empty_n;
    assign fifo_intf_2552.wr_en = AESL_inst_myproject.layer3_out_1199_U.if_write & AESL_inst_myproject.layer3_out_1199_U.if_full_n;
    assign fifo_intf_2552.fifo_rd_block = 0;
    assign fifo_intf_2552.fifo_wr_block = 0;
    assign fifo_intf_2552.finish = finish;
    csv_file_dump fifo_csv_dumper_2552;
    csv_file_dump cstatus_csv_dumper_2552;
    df_fifo_monitor fifo_monitor_2552;
    df_fifo_intf fifo_intf_2553(clock,reset);
    assign fifo_intf_2553.rd_en = AESL_inst_myproject.layer3_out_1200_U.if_read & AESL_inst_myproject.layer3_out_1200_U.if_empty_n;
    assign fifo_intf_2553.wr_en = AESL_inst_myproject.layer3_out_1200_U.if_write & AESL_inst_myproject.layer3_out_1200_U.if_full_n;
    assign fifo_intf_2553.fifo_rd_block = 0;
    assign fifo_intf_2553.fifo_wr_block = 0;
    assign fifo_intf_2553.finish = finish;
    csv_file_dump fifo_csv_dumper_2553;
    csv_file_dump cstatus_csv_dumper_2553;
    df_fifo_monitor fifo_monitor_2553;
    df_fifo_intf fifo_intf_2554(clock,reset);
    assign fifo_intf_2554.rd_en = AESL_inst_myproject.layer3_out_1201_U.if_read & AESL_inst_myproject.layer3_out_1201_U.if_empty_n;
    assign fifo_intf_2554.wr_en = AESL_inst_myproject.layer3_out_1201_U.if_write & AESL_inst_myproject.layer3_out_1201_U.if_full_n;
    assign fifo_intf_2554.fifo_rd_block = 0;
    assign fifo_intf_2554.fifo_wr_block = 0;
    assign fifo_intf_2554.finish = finish;
    csv_file_dump fifo_csv_dumper_2554;
    csv_file_dump cstatus_csv_dumper_2554;
    df_fifo_monitor fifo_monitor_2554;
    df_fifo_intf fifo_intf_2555(clock,reset);
    assign fifo_intf_2555.rd_en = AESL_inst_myproject.layer3_out_1202_U.if_read & AESL_inst_myproject.layer3_out_1202_U.if_empty_n;
    assign fifo_intf_2555.wr_en = AESL_inst_myproject.layer3_out_1202_U.if_write & AESL_inst_myproject.layer3_out_1202_U.if_full_n;
    assign fifo_intf_2555.fifo_rd_block = 0;
    assign fifo_intf_2555.fifo_wr_block = 0;
    assign fifo_intf_2555.finish = finish;
    csv_file_dump fifo_csv_dumper_2555;
    csv_file_dump cstatus_csv_dumper_2555;
    df_fifo_monitor fifo_monitor_2555;
    df_fifo_intf fifo_intf_2556(clock,reset);
    assign fifo_intf_2556.rd_en = AESL_inst_myproject.layer3_out_1203_U.if_read & AESL_inst_myproject.layer3_out_1203_U.if_empty_n;
    assign fifo_intf_2556.wr_en = AESL_inst_myproject.layer3_out_1203_U.if_write & AESL_inst_myproject.layer3_out_1203_U.if_full_n;
    assign fifo_intf_2556.fifo_rd_block = 0;
    assign fifo_intf_2556.fifo_wr_block = 0;
    assign fifo_intf_2556.finish = finish;
    csv_file_dump fifo_csv_dumper_2556;
    csv_file_dump cstatus_csv_dumper_2556;
    df_fifo_monitor fifo_monitor_2556;
    df_fifo_intf fifo_intf_2557(clock,reset);
    assign fifo_intf_2557.rd_en = AESL_inst_myproject.layer3_out_1204_U.if_read & AESL_inst_myproject.layer3_out_1204_U.if_empty_n;
    assign fifo_intf_2557.wr_en = AESL_inst_myproject.layer3_out_1204_U.if_write & AESL_inst_myproject.layer3_out_1204_U.if_full_n;
    assign fifo_intf_2557.fifo_rd_block = 0;
    assign fifo_intf_2557.fifo_wr_block = 0;
    assign fifo_intf_2557.finish = finish;
    csv_file_dump fifo_csv_dumper_2557;
    csv_file_dump cstatus_csv_dumper_2557;
    df_fifo_monitor fifo_monitor_2557;
    df_fifo_intf fifo_intf_2558(clock,reset);
    assign fifo_intf_2558.rd_en = AESL_inst_myproject.layer3_out_1205_U.if_read & AESL_inst_myproject.layer3_out_1205_U.if_empty_n;
    assign fifo_intf_2558.wr_en = AESL_inst_myproject.layer3_out_1205_U.if_write & AESL_inst_myproject.layer3_out_1205_U.if_full_n;
    assign fifo_intf_2558.fifo_rd_block = 0;
    assign fifo_intf_2558.fifo_wr_block = 0;
    assign fifo_intf_2558.finish = finish;
    csv_file_dump fifo_csv_dumper_2558;
    csv_file_dump cstatus_csv_dumper_2558;
    df_fifo_monitor fifo_monitor_2558;
    df_fifo_intf fifo_intf_2559(clock,reset);
    assign fifo_intf_2559.rd_en = AESL_inst_myproject.layer3_out_1206_U.if_read & AESL_inst_myproject.layer3_out_1206_U.if_empty_n;
    assign fifo_intf_2559.wr_en = AESL_inst_myproject.layer3_out_1206_U.if_write & AESL_inst_myproject.layer3_out_1206_U.if_full_n;
    assign fifo_intf_2559.fifo_rd_block = 0;
    assign fifo_intf_2559.fifo_wr_block = 0;
    assign fifo_intf_2559.finish = finish;
    csv_file_dump fifo_csv_dumper_2559;
    csv_file_dump cstatus_csv_dumper_2559;
    df_fifo_monitor fifo_monitor_2559;
    df_fifo_intf fifo_intf_2560(clock,reset);
    assign fifo_intf_2560.rd_en = AESL_inst_myproject.layer3_out_1207_U.if_read & AESL_inst_myproject.layer3_out_1207_U.if_empty_n;
    assign fifo_intf_2560.wr_en = AESL_inst_myproject.layer3_out_1207_U.if_write & AESL_inst_myproject.layer3_out_1207_U.if_full_n;
    assign fifo_intf_2560.fifo_rd_block = 0;
    assign fifo_intf_2560.fifo_wr_block = 0;
    assign fifo_intf_2560.finish = finish;
    csv_file_dump fifo_csv_dumper_2560;
    csv_file_dump cstatus_csv_dumper_2560;
    df_fifo_monitor fifo_monitor_2560;
    df_fifo_intf fifo_intf_2561(clock,reset);
    assign fifo_intf_2561.rd_en = AESL_inst_myproject.layer3_out_1208_U.if_read & AESL_inst_myproject.layer3_out_1208_U.if_empty_n;
    assign fifo_intf_2561.wr_en = AESL_inst_myproject.layer3_out_1208_U.if_write & AESL_inst_myproject.layer3_out_1208_U.if_full_n;
    assign fifo_intf_2561.fifo_rd_block = 0;
    assign fifo_intf_2561.fifo_wr_block = 0;
    assign fifo_intf_2561.finish = finish;
    csv_file_dump fifo_csv_dumper_2561;
    csv_file_dump cstatus_csv_dumper_2561;
    df_fifo_monitor fifo_monitor_2561;
    df_fifo_intf fifo_intf_2562(clock,reset);
    assign fifo_intf_2562.rd_en = AESL_inst_myproject.layer3_out_1209_U.if_read & AESL_inst_myproject.layer3_out_1209_U.if_empty_n;
    assign fifo_intf_2562.wr_en = AESL_inst_myproject.layer3_out_1209_U.if_write & AESL_inst_myproject.layer3_out_1209_U.if_full_n;
    assign fifo_intf_2562.fifo_rd_block = 0;
    assign fifo_intf_2562.fifo_wr_block = 0;
    assign fifo_intf_2562.finish = finish;
    csv_file_dump fifo_csv_dumper_2562;
    csv_file_dump cstatus_csv_dumper_2562;
    df_fifo_monitor fifo_monitor_2562;
    df_fifo_intf fifo_intf_2563(clock,reset);
    assign fifo_intf_2563.rd_en = AESL_inst_myproject.layer3_out_1210_U.if_read & AESL_inst_myproject.layer3_out_1210_U.if_empty_n;
    assign fifo_intf_2563.wr_en = AESL_inst_myproject.layer3_out_1210_U.if_write & AESL_inst_myproject.layer3_out_1210_U.if_full_n;
    assign fifo_intf_2563.fifo_rd_block = 0;
    assign fifo_intf_2563.fifo_wr_block = 0;
    assign fifo_intf_2563.finish = finish;
    csv_file_dump fifo_csv_dumper_2563;
    csv_file_dump cstatus_csv_dumper_2563;
    df_fifo_monitor fifo_monitor_2563;
    df_fifo_intf fifo_intf_2564(clock,reset);
    assign fifo_intf_2564.rd_en = AESL_inst_myproject.layer3_out_1211_U.if_read & AESL_inst_myproject.layer3_out_1211_U.if_empty_n;
    assign fifo_intf_2564.wr_en = AESL_inst_myproject.layer3_out_1211_U.if_write & AESL_inst_myproject.layer3_out_1211_U.if_full_n;
    assign fifo_intf_2564.fifo_rd_block = 0;
    assign fifo_intf_2564.fifo_wr_block = 0;
    assign fifo_intf_2564.finish = finish;
    csv_file_dump fifo_csv_dumper_2564;
    csv_file_dump cstatus_csv_dumper_2564;
    df_fifo_monitor fifo_monitor_2564;
    df_fifo_intf fifo_intf_2565(clock,reset);
    assign fifo_intf_2565.rd_en = AESL_inst_myproject.layer3_out_1212_U.if_read & AESL_inst_myproject.layer3_out_1212_U.if_empty_n;
    assign fifo_intf_2565.wr_en = AESL_inst_myproject.layer3_out_1212_U.if_write & AESL_inst_myproject.layer3_out_1212_U.if_full_n;
    assign fifo_intf_2565.fifo_rd_block = 0;
    assign fifo_intf_2565.fifo_wr_block = 0;
    assign fifo_intf_2565.finish = finish;
    csv_file_dump fifo_csv_dumper_2565;
    csv_file_dump cstatus_csv_dumper_2565;
    df_fifo_monitor fifo_monitor_2565;
    df_fifo_intf fifo_intf_2566(clock,reset);
    assign fifo_intf_2566.rd_en = AESL_inst_myproject.layer3_out_1213_U.if_read & AESL_inst_myproject.layer3_out_1213_U.if_empty_n;
    assign fifo_intf_2566.wr_en = AESL_inst_myproject.layer3_out_1213_U.if_write & AESL_inst_myproject.layer3_out_1213_U.if_full_n;
    assign fifo_intf_2566.fifo_rd_block = 0;
    assign fifo_intf_2566.fifo_wr_block = 0;
    assign fifo_intf_2566.finish = finish;
    csv_file_dump fifo_csv_dumper_2566;
    csv_file_dump cstatus_csv_dumper_2566;
    df_fifo_monitor fifo_monitor_2566;
    df_fifo_intf fifo_intf_2567(clock,reset);
    assign fifo_intf_2567.rd_en = AESL_inst_myproject.layer3_out_1214_U.if_read & AESL_inst_myproject.layer3_out_1214_U.if_empty_n;
    assign fifo_intf_2567.wr_en = AESL_inst_myproject.layer3_out_1214_U.if_write & AESL_inst_myproject.layer3_out_1214_U.if_full_n;
    assign fifo_intf_2567.fifo_rd_block = 0;
    assign fifo_intf_2567.fifo_wr_block = 0;
    assign fifo_intf_2567.finish = finish;
    csv_file_dump fifo_csv_dumper_2567;
    csv_file_dump cstatus_csv_dumper_2567;
    df_fifo_monitor fifo_monitor_2567;
    df_fifo_intf fifo_intf_2568(clock,reset);
    assign fifo_intf_2568.rd_en = AESL_inst_myproject.layer3_out_1215_U.if_read & AESL_inst_myproject.layer3_out_1215_U.if_empty_n;
    assign fifo_intf_2568.wr_en = AESL_inst_myproject.layer3_out_1215_U.if_write & AESL_inst_myproject.layer3_out_1215_U.if_full_n;
    assign fifo_intf_2568.fifo_rd_block = 0;
    assign fifo_intf_2568.fifo_wr_block = 0;
    assign fifo_intf_2568.finish = finish;
    csv_file_dump fifo_csv_dumper_2568;
    csv_file_dump cstatus_csv_dumper_2568;
    df_fifo_monitor fifo_monitor_2568;
    df_fifo_intf fifo_intf_2569(clock,reset);
    assign fifo_intf_2569.rd_en = AESL_inst_myproject.layer3_out_1216_U.if_read & AESL_inst_myproject.layer3_out_1216_U.if_empty_n;
    assign fifo_intf_2569.wr_en = AESL_inst_myproject.layer3_out_1216_U.if_write & AESL_inst_myproject.layer3_out_1216_U.if_full_n;
    assign fifo_intf_2569.fifo_rd_block = 0;
    assign fifo_intf_2569.fifo_wr_block = 0;
    assign fifo_intf_2569.finish = finish;
    csv_file_dump fifo_csv_dumper_2569;
    csv_file_dump cstatus_csv_dumper_2569;
    df_fifo_monitor fifo_monitor_2569;
    df_fifo_intf fifo_intf_2570(clock,reset);
    assign fifo_intf_2570.rd_en = AESL_inst_myproject.layer3_out_1217_U.if_read & AESL_inst_myproject.layer3_out_1217_U.if_empty_n;
    assign fifo_intf_2570.wr_en = AESL_inst_myproject.layer3_out_1217_U.if_write & AESL_inst_myproject.layer3_out_1217_U.if_full_n;
    assign fifo_intf_2570.fifo_rd_block = 0;
    assign fifo_intf_2570.fifo_wr_block = 0;
    assign fifo_intf_2570.finish = finish;
    csv_file_dump fifo_csv_dumper_2570;
    csv_file_dump cstatus_csv_dumper_2570;
    df_fifo_monitor fifo_monitor_2570;
    df_fifo_intf fifo_intf_2571(clock,reset);
    assign fifo_intf_2571.rd_en = AESL_inst_myproject.layer3_out_1218_U.if_read & AESL_inst_myproject.layer3_out_1218_U.if_empty_n;
    assign fifo_intf_2571.wr_en = AESL_inst_myproject.layer3_out_1218_U.if_write & AESL_inst_myproject.layer3_out_1218_U.if_full_n;
    assign fifo_intf_2571.fifo_rd_block = 0;
    assign fifo_intf_2571.fifo_wr_block = 0;
    assign fifo_intf_2571.finish = finish;
    csv_file_dump fifo_csv_dumper_2571;
    csv_file_dump cstatus_csv_dumper_2571;
    df_fifo_monitor fifo_monitor_2571;
    df_fifo_intf fifo_intf_2572(clock,reset);
    assign fifo_intf_2572.rd_en = AESL_inst_myproject.layer3_out_1219_U.if_read & AESL_inst_myproject.layer3_out_1219_U.if_empty_n;
    assign fifo_intf_2572.wr_en = AESL_inst_myproject.layer3_out_1219_U.if_write & AESL_inst_myproject.layer3_out_1219_U.if_full_n;
    assign fifo_intf_2572.fifo_rd_block = 0;
    assign fifo_intf_2572.fifo_wr_block = 0;
    assign fifo_intf_2572.finish = finish;
    csv_file_dump fifo_csv_dumper_2572;
    csv_file_dump cstatus_csv_dumper_2572;
    df_fifo_monitor fifo_monitor_2572;
    df_fifo_intf fifo_intf_2573(clock,reset);
    assign fifo_intf_2573.rd_en = AESL_inst_myproject.layer3_out_1220_U.if_read & AESL_inst_myproject.layer3_out_1220_U.if_empty_n;
    assign fifo_intf_2573.wr_en = AESL_inst_myproject.layer3_out_1220_U.if_write & AESL_inst_myproject.layer3_out_1220_U.if_full_n;
    assign fifo_intf_2573.fifo_rd_block = 0;
    assign fifo_intf_2573.fifo_wr_block = 0;
    assign fifo_intf_2573.finish = finish;
    csv_file_dump fifo_csv_dumper_2573;
    csv_file_dump cstatus_csv_dumper_2573;
    df_fifo_monitor fifo_monitor_2573;
    df_fifo_intf fifo_intf_2574(clock,reset);
    assign fifo_intf_2574.rd_en = AESL_inst_myproject.layer3_out_1221_U.if_read & AESL_inst_myproject.layer3_out_1221_U.if_empty_n;
    assign fifo_intf_2574.wr_en = AESL_inst_myproject.layer3_out_1221_U.if_write & AESL_inst_myproject.layer3_out_1221_U.if_full_n;
    assign fifo_intf_2574.fifo_rd_block = 0;
    assign fifo_intf_2574.fifo_wr_block = 0;
    assign fifo_intf_2574.finish = finish;
    csv_file_dump fifo_csv_dumper_2574;
    csv_file_dump cstatus_csv_dumper_2574;
    df_fifo_monitor fifo_monitor_2574;
    df_fifo_intf fifo_intf_2575(clock,reset);
    assign fifo_intf_2575.rd_en = AESL_inst_myproject.layer3_out_1222_U.if_read & AESL_inst_myproject.layer3_out_1222_U.if_empty_n;
    assign fifo_intf_2575.wr_en = AESL_inst_myproject.layer3_out_1222_U.if_write & AESL_inst_myproject.layer3_out_1222_U.if_full_n;
    assign fifo_intf_2575.fifo_rd_block = 0;
    assign fifo_intf_2575.fifo_wr_block = 0;
    assign fifo_intf_2575.finish = finish;
    csv_file_dump fifo_csv_dumper_2575;
    csv_file_dump cstatus_csv_dumper_2575;
    df_fifo_monitor fifo_monitor_2575;
    df_fifo_intf fifo_intf_2576(clock,reset);
    assign fifo_intf_2576.rd_en = AESL_inst_myproject.layer3_out_1223_U.if_read & AESL_inst_myproject.layer3_out_1223_U.if_empty_n;
    assign fifo_intf_2576.wr_en = AESL_inst_myproject.layer3_out_1223_U.if_write & AESL_inst_myproject.layer3_out_1223_U.if_full_n;
    assign fifo_intf_2576.fifo_rd_block = 0;
    assign fifo_intf_2576.fifo_wr_block = 0;
    assign fifo_intf_2576.finish = finish;
    csv_file_dump fifo_csv_dumper_2576;
    csv_file_dump cstatus_csv_dumper_2576;
    df_fifo_monitor fifo_monitor_2576;
    df_fifo_intf fifo_intf_2577(clock,reset);
    assign fifo_intf_2577.rd_en = AESL_inst_myproject.layer3_out_1224_U.if_read & AESL_inst_myproject.layer3_out_1224_U.if_empty_n;
    assign fifo_intf_2577.wr_en = AESL_inst_myproject.layer3_out_1224_U.if_write & AESL_inst_myproject.layer3_out_1224_U.if_full_n;
    assign fifo_intf_2577.fifo_rd_block = 0;
    assign fifo_intf_2577.fifo_wr_block = 0;
    assign fifo_intf_2577.finish = finish;
    csv_file_dump fifo_csv_dumper_2577;
    csv_file_dump cstatus_csv_dumper_2577;
    df_fifo_monitor fifo_monitor_2577;
    df_fifo_intf fifo_intf_2578(clock,reset);
    assign fifo_intf_2578.rd_en = AESL_inst_myproject.layer3_out_1225_U.if_read & AESL_inst_myproject.layer3_out_1225_U.if_empty_n;
    assign fifo_intf_2578.wr_en = AESL_inst_myproject.layer3_out_1225_U.if_write & AESL_inst_myproject.layer3_out_1225_U.if_full_n;
    assign fifo_intf_2578.fifo_rd_block = 0;
    assign fifo_intf_2578.fifo_wr_block = 0;
    assign fifo_intf_2578.finish = finish;
    csv_file_dump fifo_csv_dumper_2578;
    csv_file_dump cstatus_csv_dumper_2578;
    df_fifo_monitor fifo_monitor_2578;
    df_fifo_intf fifo_intf_2579(clock,reset);
    assign fifo_intf_2579.rd_en = AESL_inst_myproject.layer3_out_1226_U.if_read & AESL_inst_myproject.layer3_out_1226_U.if_empty_n;
    assign fifo_intf_2579.wr_en = AESL_inst_myproject.layer3_out_1226_U.if_write & AESL_inst_myproject.layer3_out_1226_U.if_full_n;
    assign fifo_intf_2579.fifo_rd_block = 0;
    assign fifo_intf_2579.fifo_wr_block = 0;
    assign fifo_intf_2579.finish = finish;
    csv_file_dump fifo_csv_dumper_2579;
    csv_file_dump cstatus_csv_dumper_2579;
    df_fifo_monitor fifo_monitor_2579;
    df_fifo_intf fifo_intf_2580(clock,reset);
    assign fifo_intf_2580.rd_en = AESL_inst_myproject.layer3_out_1227_U.if_read & AESL_inst_myproject.layer3_out_1227_U.if_empty_n;
    assign fifo_intf_2580.wr_en = AESL_inst_myproject.layer3_out_1227_U.if_write & AESL_inst_myproject.layer3_out_1227_U.if_full_n;
    assign fifo_intf_2580.fifo_rd_block = 0;
    assign fifo_intf_2580.fifo_wr_block = 0;
    assign fifo_intf_2580.finish = finish;
    csv_file_dump fifo_csv_dumper_2580;
    csv_file_dump cstatus_csv_dumper_2580;
    df_fifo_monitor fifo_monitor_2580;
    df_fifo_intf fifo_intf_2581(clock,reset);
    assign fifo_intf_2581.rd_en = AESL_inst_myproject.layer3_out_1228_U.if_read & AESL_inst_myproject.layer3_out_1228_U.if_empty_n;
    assign fifo_intf_2581.wr_en = AESL_inst_myproject.layer3_out_1228_U.if_write & AESL_inst_myproject.layer3_out_1228_U.if_full_n;
    assign fifo_intf_2581.fifo_rd_block = 0;
    assign fifo_intf_2581.fifo_wr_block = 0;
    assign fifo_intf_2581.finish = finish;
    csv_file_dump fifo_csv_dumper_2581;
    csv_file_dump cstatus_csv_dumper_2581;
    df_fifo_monitor fifo_monitor_2581;
    df_fifo_intf fifo_intf_2582(clock,reset);
    assign fifo_intf_2582.rd_en = AESL_inst_myproject.layer3_out_1229_U.if_read & AESL_inst_myproject.layer3_out_1229_U.if_empty_n;
    assign fifo_intf_2582.wr_en = AESL_inst_myproject.layer3_out_1229_U.if_write & AESL_inst_myproject.layer3_out_1229_U.if_full_n;
    assign fifo_intf_2582.fifo_rd_block = 0;
    assign fifo_intf_2582.fifo_wr_block = 0;
    assign fifo_intf_2582.finish = finish;
    csv_file_dump fifo_csv_dumper_2582;
    csv_file_dump cstatus_csv_dumper_2582;
    df_fifo_monitor fifo_monitor_2582;
    df_fifo_intf fifo_intf_2583(clock,reset);
    assign fifo_intf_2583.rd_en = AESL_inst_myproject.layer3_out_1230_U.if_read & AESL_inst_myproject.layer3_out_1230_U.if_empty_n;
    assign fifo_intf_2583.wr_en = AESL_inst_myproject.layer3_out_1230_U.if_write & AESL_inst_myproject.layer3_out_1230_U.if_full_n;
    assign fifo_intf_2583.fifo_rd_block = 0;
    assign fifo_intf_2583.fifo_wr_block = 0;
    assign fifo_intf_2583.finish = finish;
    csv_file_dump fifo_csv_dumper_2583;
    csv_file_dump cstatus_csv_dumper_2583;
    df_fifo_monitor fifo_monitor_2583;
    df_fifo_intf fifo_intf_2584(clock,reset);
    assign fifo_intf_2584.rd_en = AESL_inst_myproject.layer3_out_1231_U.if_read & AESL_inst_myproject.layer3_out_1231_U.if_empty_n;
    assign fifo_intf_2584.wr_en = AESL_inst_myproject.layer3_out_1231_U.if_write & AESL_inst_myproject.layer3_out_1231_U.if_full_n;
    assign fifo_intf_2584.fifo_rd_block = 0;
    assign fifo_intf_2584.fifo_wr_block = 0;
    assign fifo_intf_2584.finish = finish;
    csv_file_dump fifo_csv_dumper_2584;
    csv_file_dump cstatus_csv_dumper_2584;
    df_fifo_monitor fifo_monitor_2584;
    df_fifo_intf fifo_intf_2585(clock,reset);
    assign fifo_intf_2585.rd_en = AESL_inst_myproject.layer3_out_1232_U.if_read & AESL_inst_myproject.layer3_out_1232_U.if_empty_n;
    assign fifo_intf_2585.wr_en = AESL_inst_myproject.layer3_out_1232_U.if_write & AESL_inst_myproject.layer3_out_1232_U.if_full_n;
    assign fifo_intf_2585.fifo_rd_block = 0;
    assign fifo_intf_2585.fifo_wr_block = 0;
    assign fifo_intf_2585.finish = finish;
    csv_file_dump fifo_csv_dumper_2585;
    csv_file_dump cstatus_csv_dumper_2585;
    df_fifo_monitor fifo_monitor_2585;
    df_fifo_intf fifo_intf_2586(clock,reset);
    assign fifo_intf_2586.rd_en = AESL_inst_myproject.layer3_out_1233_U.if_read & AESL_inst_myproject.layer3_out_1233_U.if_empty_n;
    assign fifo_intf_2586.wr_en = AESL_inst_myproject.layer3_out_1233_U.if_write & AESL_inst_myproject.layer3_out_1233_U.if_full_n;
    assign fifo_intf_2586.fifo_rd_block = 0;
    assign fifo_intf_2586.fifo_wr_block = 0;
    assign fifo_intf_2586.finish = finish;
    csv_file_dump fifo_csv_dumper_2586;
    csv_file_dump cstatus_csv_dumper_2586;
    df_fifo_monitor fifo_monitor_2586;
    df_fifo_intf fifo_intf_2587(clock,reset);
    assign fifo_intf_2587.rd_en = AESL_inst_myproject.layer3_out_1234_U.if_read & AESL_inst_myproject.layer3_out_1234_U.if_empty_n;
    assign fifo_intf_2587.wr_en = AESL_inst_myproject.layer3_out_1234_U.if_write & AESL_inst_myproject.layer3_out_1234_U.if_full_n;
    assign fifo_intf_2587.fifo_rd_block = 0;
    assign fifo_intf_2587.fifo_wr_block = 0;
    assign fifo_intf_2587.finish = finish;
    csv_file_dump fifo_csv_dumper_2587;
    csv_file_dump cstatus_csv_dumper_2587;
    df_fifo_monitor fifo_monitor_2587;
    df_fifo_intf fifo_intf_2588(clock,reset);
    assign fifo_intf_2588.rd_en = AESL_inst_myproject.layer3_out_1235_U.if_read & AESL_inst_myproject.layer3_out_1235_U.if_empty_n;
    assign fifo_intf_2588.wr_en = AESL_inst_myproject.layer3_out_1235_U.if_write & AESL_inst_myproject.layer3_out_1235_U.if_full_n;
    assign fifo_intf_2588.fifo_rd_block = 0;
    assign fifo_intf_2588.fifo_wr_block = 0;
    assign fifo_intf_2588.finish = finish;
    csv_file_dump fifo_csv_dumper_2588;
    csv_file_dump cstatus_csv_dumper_2588;
    df_fifo_monitor fifo_monitor_2588;
    df_fifo_intf fifo_intf_2589(clock,reset);
    assign fifo_intf_2589.rd_en = AESL_inst_myproject.layer3_out_1236_U.if_read & AESL_inst_myproject.layer3_out_1236_U.if_empty_n;
    assign fifo_intf_2589.wr_en = AESL_inst_myproject.layer3_out_1236_U.if_write & AESL_inst_myproject.layer3_out_1236_U.if_full_n;
    assign fifo_intf_2589.fifo_rd_block = 0;
    assign fifo_intf_2589.fifo_wr_block = 0;
    assign fifo_intf_2589.finish = finish;
    csv_file_dump fifo_csv_dumper_2589;
    csv_file_dump cstatus_csv_dumper_2589;
    df_fifo_monitor fifo_monitor_2589;
    df_fifo_intf fifo_intf_2590(clock,reset);
    assign fifo_intf_2590.rd_en = AESL_inst_myproject.layer3_out_1237_U.if_read & AESL_inst_myproject.layer3_out_1237_U.if_empty_n;
    assign fifo_intf_2590.wr_en = AESL_inst_myproject.layer3_out_1237_U.if_write & AESL_inst_myproject.layer3_out_1237_U.if_full_n;
    assign fifo_intf_2590.fifo_rd_block = 0;
    assign fifo_intf_2590.fifo_wr_block = 0;
    assign fifo_intf_2590.finish = finish;
    csv_file_dump fifo_csv_dumper_2590;
    csv_file_dump cstatus_csv_dumper_2590;
    df_fifo_monitor fifo_monitor_2590;
    df_fifo_intf fifo_intf_2591(clock,reset);
    assign fifo_intf_2591.rd_en = AESL_inst_myproject.layer3_out_1238_U.if_read & AESL_inst_myproject.layer3_out_1238_U.if_empty_n;
    assign fifo_intf_2591.wr_en = AESL_inst_myproject.layer3_out_1238_U.if_write & AESL_inst_myproject.layer3_out_1238_U.if_full_n;
    assign fifo_intf_2591.fifo_rd_block = 0;
    assign fifo_intf_2591.fifo_wr_block = 0;
    assign fifo_intf_2591.finish = finish;
    csv_file_dump fifo_csv_dumper_2591;
    csv_file_dump cstatus_csv_dumper_2591;
    df_fifo_monitor fifo_monitor_2591;
    df_fifo_intf fifo_intf_2592(clock,reset);
    assign fifo_intf_2592.rd_en = AESL_inst_myproject.layer3_out_1239_U.if_read & AESL_inst_myproject.layer3_out_1239_U.if_empty_n;
    assign fifo_intf_2592.wr_en = AESL_inst_myproject.layer3_out_1239_U.if_write & AESL_inst_myproject.layer3_out_1239_U.if_full_n;
    assign fifo_intf_2592.fifo_rd_block = 0;
    assign fifo_intf_2592.fifo_wr_block = 0;
    assign fifo_intf_2592.finish = finish;
    csv_file_dump fifo_csv_dumper_2592;
    csv_file_dump cstatus_csv_dumper_2592;
    df_fifo_monitor fifo_monitor_2592;
    df_fifo_intf fifo_intf_2593(clock,reset);
    assign fifo_intf_2593.rd_en = AESL_inst_myproject.layer3_out_1240_U.if_read & AESL_inst_myproject.layer3_out_1240_U.if_empty_n;
    assign fifo_intf_2593.wr_en = AESL_inst_myproject.layer3_out_1240_U.if_write & AESL_inst_myproject.layer3_out_1240_U.if_full_n;
    assign fifo_intf_2593.fifo_rd_block = 0;
    assign fifo_intf_2593.fifo_wr_block = 0;
    assign fifo_intf_2593.finish = finish;
    csv_file_dump fifo_csv_dumper_2593;
    csv_file_dump cstatus_csv_dumper_2593;
    df_fifo_monitor fifo_monitor_2593;
    df_fifo_intf fifo_intf_2594(clock,reset);
    assign fifo_intf_2594.rd_en = AESL_inst_myproject.layer3_out_1241_U.if_read & AESL_inst_myproject.layer3_out_1241_U.if_empty_n;
    assign fifo_intf_2594.wr_en = AESL_inst_myproject.layer3_out_1241_U.if_write & AESL_inst_myproject.layer3_out_1241_U.if_full_n;
    assign fifo_intf_2594.fifo_rd_block = 0;
    assign fifo_intf_2594.fifo_wr_block = 0;
    assign fifo_intf_2594.finish = finish;
    csv_file_dump fifo_csv_dumper_2594;
    csv_file_dump cstatus_csv_dumper_2594;
    df_fifo_monitor fifo_monitor_2594;
    df_fifo_intf fifo_intf_2595(clock,reset);
    assign fifo_intf_2595.rd_en = AESL_inst_myproject.layer3_out_1242_U.if_read & AESL_inst_myproject.layer3_out_1242_U.if_empty_n;
    assign fifo_intf_2595.wr_en = AESL_inst_myproject.layer3_out_1242_U.if_write & AESL_inst_myproject.layer3_out_1242_U.if_full_n;
    assign fifo_intf_2595.fifo_rd_block = 0;
    assign fifo_intf_2595.fifo_wr_block = 0;
    assign fifo_intf_2595.finish = finish;
    csv_file_dump fifo_csv_dumper_2595;
    csv_file_dump cstatus_csv_dumper_2595;
    df_fifo_monitor fifo_monitor_2595;
    df_fifo_intf fifo_intf_2596(clock,reset);
    assign fifo_intf_2596.rd_en = AESL_inst_myproject.layer3_out_1243_U.if_read & AESL_inst_myproject.layer3_out_1243_U.if_empty_n;
    assign fifo_intf_2596.wr_en = AESL_inst_myproject.layer3_out_1243_U.if_write & AESL_inst_myproject.layer3_out_1243_U.if_full_n;
    assign fifo_intf_2596.fifo_rd_block = 0;
    assign fifo_intf_2596.fifo_wr_block = 0;
    assign fifo_intf_2596.finish = finish;
    csv_file_dump fifo_csv_dumper_2596;
    csv_file_dump cstatus_csv_dumper_2596;
    df_fifo_monitor fifo_monitor_2596;
    df_fifo_intf fifo_intf_2597(clock,reset);
    assign fifo_intf_2597.rd_en = AESL_inst_myproject.layer3_out_1244_U.if_read & AESL_inst_myproject.layer3_out_1244_U.if_empty_n;
    assign fifo_intf_2597.wr_en = AESL_inst_myproject.layer3_out_1244_U.if_write & AESL_inst_myproject.layer3_out_1244_U.if_full_n;
    assign fifo_intf_2597.fifo_rd_block = 0;
    assign fifo_intf_2597.fifo_wr_block = 0;
    assign fifo_intf_2597.finish = finish;
    csv_file_dump fifo_csv_dumper_2597;
    csv_file_dump cstatus_csv_dumper_2597;
    df_fifo_monitor fifo_monitor_2597;
    df_fifo_intf fifo_intf_2598(clock,reset);
    assign fifo_intf_2598.rd_en = AESL_inst_myproject.layer3_out_1245_U.if_read & AESL_inst_myproject.layer3_out_1245_U.if_empty_n;
    assign fifo_intf_2598.wr_en = AESL_inst_myproject.layer3_out_1245_U.if_write & AESL_inst_myproject.layer3_out_1245_U.if_full_n;
    assign fifo_intf_2598.fifo_rd_block = 0;
    assign fifo_intf_2598.fifo_wr_block = 0;
    assign fifo_intf_2598.finish = finish;
    csv_file_dump fifo_csv_dumper_2598;
    csv_file_dump cstatus_csv_dumper_2598;
    df_fifo_monitor fifo_monitor_2598;
    df_fifo_intf fifo_intf_2599(clock,reset);
    assign fifo_intf_2599.rd_en = AESL_inst_myproject.layer3_out_1246_U.if_read & AESL_inst_myproject.layer3_out_1246_U.if_empty_n;
    assign fifo_intf_2599.wr_en = AESL_inst_myproject.layer3_out_1246_U.if_write & AESL_inst_myproject.layer3_out_1246_U.if_full_n;
    assign fifo_intf_2599.fifo_rd_block = 0;
    assign fifo_intf_2599.fifo_wr_block = 0;
    assign fifo_intf_2599.finish = finish;
    csv_file_dump fifo_csv_dumper_2599;
    csv_file_dump cstatus_csv_dumper_2599;
    df_fifo_monitor fifo_monitor_2599;
    df_fifo_intf fifo_intf_2600(clock,reset);
    assign fifo_intf_2600.rd_en = AESL_inst_myproject.layer3_out_1247_U.if_read & AESL_inst_myproject.layer3_out_1247_U.if_empty_n;
    assign fifo_intf_2600.wr_en = AESL_inst_myproject.layer3_out_1247_U.if_write & AESL_inst_myproject.layer3_out_1247_U.if_full_n;
    assign fifo_intf_2600.fifo_rd_block = 0;
    assign fifo_intf_2600.fifo_wr_block = 0;
    assign fifo_intf_2600.finish = finish;
    csv_file_dump fifo_csv_dumper_2600;
    csv_file_dump cstatus_csv_dumper_2600;
    df_fifo_monitor fifo_monitor_2600;
    df_fifo_intf fifo_intf_2601(clock,reset);
    assign fifo_intf_2601.rd_en = AESL_inst_myproject.layer3_out_1248_U.if_read & AESL_inst_myproject.layer3_out_1248_U.if_empty_n;
    assign fifo_intf_2601.wr_en = AESL_inst_myproject.layer3_out_1248_U.if_write & AESL_inst_myproject.layer3_out_1248_U.if_full_n;
    assign fifo_intf_2601.fifo_rd_block = 0;
    assign fifo_intf_2601.fifo_wr_block = 0;
    assign fifo_intf_2601.finish = finish;
    csv_file_dump fifo_csv_dumper_2601;
    csv_file_dump cstatus_csv_dumper_2601;
    df_fifo_monitor fifo_monitor_2601;
    df_fifo_intf fifo_intf_2602(clock,reset);
    assign fifo_intf_2602.rd_en = AESL_inst_myproject.layer3_out_1249_U.if_read & AESL_inst_myproject.layer3_out_1249_U.if_empty_n;
    assign fifo_intf_2602.wr_en = AESL_inst_myproject.layer3_out_1249_U.if_write & AESL_inst_myproject.layer3_out_1249_U.if_full_n;
    assign fifo_intf_2602.fifo_rd_block = 0;
    assign fifo_intf_2602.fifo_wr_block = 0;
    assign fifo_intf_2602.finish = finish;
    csv_file_dump fifo_csv_dumper_2602;
    csv_file_dump cstatus_csv_dumper_2602;
    df_fifo_monitor fifo_monitor_2602;
    df_fifo_intf fifo_intf_2603(clock,reset);
    assign fifo_intf_2603.rd_en = AESL_inst_myproject.layer3_out_1250_U.if_read & AESL_inst_myproject.layer3_out_1250_U.if_empty_n;
    assign fifo_intf_2603.wr_en = AESL_inst_myproject.layer3_out_1250_U.if_write & AESL_inst_myproject.layer3_out_1250_U.if_full_n;
    assign fifo_intf_2603.fifo_rd_block = 0;
    assign fifo_intf_2603.fifo_wr_block = 0;
    assign fifo_intf_2603.finish = finish;
    csv_file_dump fifo_csv_dumper_2603;
    csv_file_dump cstatus_csv_dumper_2603;
    df_fifo_monitor fifo_monitor_2603;
    df_fifo_intf fifo_intf_2604(clock,reset);
    assign fifo_intf_2604.rd_en = AESL_inst_myproject.layer3_out_1251_U.if_read & AESL_inst_myproject.layer3_out_1251_U.if_empty_n;
    assign fifo_intf_2604.wr_en = AESL_inst_myproject.layer3_out_1251_U.if_write & AESL_inst_myproject.layer3_out_1251_U.if_full_n;
    assign fifo_intf_2604.fifo_rd_block = 0;
    assign fifo_intf_2604.fifo_wr_block = 0;
    assign fifo_intf_2604.finish = finish;
    csv_file_dump fifo_csv_dumper_2604;
    csv_file_dump cstatus_csv_dumper_2604;
    df_fifo_monitor fifo_monitor_2604;
    df_fifo_intf fifo_intf_2605(clock,reset);
    assign fifo_intf_2605.rd_en = AESL_inst_myproject.layer3_out_1252_U.if_read & AESL_inst_myproject.layer3_out_1252_U.if_empty_n;
    assign fifo_intf_2605.wr_en = AESL_inst_myproject.layer3_out_1252_U.if_write & AESL_inst_myproject.layer3_out_1252_U.if_full_n;
    assign fifo_intf_2605.fifo_rd_block = 0;
    assign fifo_intf_2605.fifo_wr_block = 0;
    assign fifo_intf_2605.finish = finish;
    csv_file_dump fifo_csv_dumper_2605;
    csv_file_dump cstatus_csv_dumper_2605;
    df_fifo_monitor fifo_monitor_2605;
    df_fifo_intf fifo_intf_2606(clock,reset);
    assign fifo_intf_2606.rd_en = AESL_inst_myproject.layer3_out_1253_U.if_read & AESL_inst_myproject.layer3_out_1253_U.if_empty_n;
    assign fifo_intf_2606.wr_en = AESL_inst_myproject.layer3_out_1253_U.if_write & AESL_inst_myproject.layer3_out_1253_U.if_full_n;
    assign fifo_intf_2606.fifo_rd_block = 0;
    assign fifo_intf_2606.fifo_wr_block = 0;
    assign fifo_intf_2606.finish = finish;
    csv_file_dump fifo_csv_dumper_2606;
    csv_file_dump cstatus_csv_dumper_2606;
    df_fifo_monitor fifo_monitor_2606;
    df_fifo_intf fifo_intf_2607(clock,reset);
    assign fifo_intf_2607.rd_en = AESL_inst_myproject.layer3_out_1254_U.if_read & AESL_inst_myproject.layer3_out_1254_U.if_empty_n;
    assign fifo_intf_2607.wr_en = AESL_inst_myproject.layer3_out_1254_U.if_write & AESL_inst_myproject.layer3_out_1254_U.if_full_n;
    assign fifo_intf_2607.fifo_rd_block = 0;
    assign fifo_intf_2607.fifo_wr_block = 0;
    assign fifo_intf_2607.finish = finish;
    csv_file_dump fifo_csv_dumper_2607;
    csv_file_dump cstatus_csv_dumper_2607;
    df_fifo_monitor fifo_monitor_2607;
    df_fifo_intf fifo_intf_2608(clock,reset);
    assign fifo_intf_2608.rd_en = AESL_inst_myproject.layer3_out_1255_U.if_read & AESL_inst_myproject.layer3_out_1255_U.if_empty_n;
    assign fifo_intf_2608.wr_en = AESL_inst_myproject.layer3_out_1255_U.if_write & AESL_inst_myproject.layer3_out_1255_U.if_full_n;
    assign fifo_intf_2608.fifo_rd_block = 0;
    assign fifo_intf_2608.fifo_wr_block = 0;
    assign fifo_intf_2608.finish = finish;
    csv_file_dump fifo_csv_dumper_2608;
    csv_file_dump cstatus_csv_dumper_2608;
    df_fifo_monitor fifo_monitor_2608;
    df_fifo_intf fifo_intf_2609(clock,reset);
    assign fifo_intf_2609.rd_en = AESL_inst_myproject.layer3_out_1256_U.if_read & AESL_inst_myproject.layer3_out_1256_U.if_empty_n;
    assign fifo_intf_2609.wr_en = AESL_inst_myproject.layer3_out_1256_U.if_write & AESL_inst_myproject.layer3_out_1256_U.if_full_n;
    assign fifo_intf_2609.fifo_rd_block = 0;
    assign fifo_intf_2609.fifo_wr_block = 0;
    assign fifo_intf_2609.finish = finish;
    csv_file_dump fifo_csv_dumper_2609;
    csv_file_dump cstatus_csv_dumper_2609;
    df_fifo_monitor fifo_monitor_2609;
    df_fifo_intf fifo_intf_2610(clock,reset);
    assign fifo_intf_2610.rd_en = AESL_inst_myproject.layer3_out_1257_U.if_read & AESL_inst_myproject.layer3_out_1257_U.if_empty_n;
    assign fifo_intf_2610.wr_en = AESL_inst_myproject.layer3_out_1257_U.if_write & AESL_inst_myproject.layer3_out_1257_U.if_full_n;
    assign fifo_intf_2610.fifo_rd_block = 0;
    assign fifo_intf_2610.fifo_wr_block = 0;
    assign fifo_intf_2610.finish = finish;
    csv_file_dump fifo_csv_dumper_2610;
    csv_file_dump cstatus_csv_dumper_2610;
    df_fifo_monitor fifo_monitor_2610;
    df_fifo_intf fifo_intf_2611(clock,reset);
    assign fifo_intf_2611.rd_en = AESL_inst_myproject.layer3_out_1258_U.if_read & AESL_inst_myproject.layer3_out_1258_U.if_empty_n;
    assign fifo_intf_2611.wr_en = AESL_inst_myproject.layer3_out_1258_U.if_write & AESL_inst_myproject.layer3_out_1258_U.if_full_n;
    assign fifo_intf_2611.fifo_rd_block = 0;
    assign fifo_intf_2611.fifo_wr_block = 0;
    assign fifo_intf_2611.finish = finish;
    csv_file_dump fifo_csv_dumper_2611;
    csv_file_dump cstatus_csv_dumper_2611;
    df_fifo_monitor fifo_monitor_2611;
    df_fifo_intf fifo_intf_2612(clock,reset);
    assign fifo_intf_2612.rd_en = AESL_inst_myproject.layer3_out_1259_U.if_read & AESL_inst_myproject.layer3_out_1259_U.if_empty_n;
    assign fifo_intf_2612.wr_en = AESL_inst_myproject.layer3_out_1259_U.if_write & AESL_inst_myproject.layer3_out_1259_U.if_full_n;
    assign fifo_intf_2612.fifo_rd_block = 0;
    assign fifo_intf_2612.fifo_wr_block = 0;
    assign fifo_intf_2612.finish = finish;
    csv_file_dump fifo_csv_dumper_2612;
    csv_file_dump cstatus_csv_dumper_2612;
    df_fifo_monitor fifo_monitor_2612;
    df_fifo_intf fifo_intf_2613(clock,reset);
    assign fifo_intf_2613.rd_en = AESL_inst_myproject.layer3_out_1260_U.if_read & AESL_inst_myproject.layer3_out_1260_U.if_empty_n;
    assign fifo_intf_2613.wr_en = AESL_inst_myproject.layer3_out_1260_U.if_write & AESL_inst_myproject.layer3_out_1260_U.if_full_n;
    assign fifo_intf_2613.fifo_rd_block = 0;
    assign fifo_intf_2613.fifo_wr_block = 0;
    assign fifo_intf_2613.finish = finish;
    csv_file_dump fifo_csv_dumper_2613;
    csv_file_dump cstatus_csv_dumper_2613;
    df_fifo_monitor fifo_monitor_2613;
    df_fifo_intf fifo_intf_2614(clock,reset);
    assign fifo_intf_2614.rd_en = AESL_inst_myproject.layer3_out_1261_U.if_read & AESL_inst_myproject.layer3_out_1261_U.if_empty_n;
    assign fifo_intf_2614.wr_en = AESL_inst_myproject.layer3_out_1261_U.if_write & AESL_inst_myproject.layer3_out_1261_U.if_full_n;
    assign fifo_intf_2614.fifo_rd_block = 0;
    assign fifo_intf_2614.fifo_wr_block = 0;
    assign fifo_intf_2614.finish = finish;
    csv_file_dump fifo_csv_dumper_2614;
    csv_file_dump cstatus_csv_dumper_2614;
    df_fifo_monitor fifo_monitor_2614;
    df_fifo_intf fifo_intf_2615(clock,reset);
    assign fifo_intf_2615.rd_en = AESL_inst_myproject.layer3_out_1262_U.if_read & AESL_inst_myproject.layer3_out_1262_U.if_empty_n;
    assign fifo_intf_2615.wr_en = AESL_inst_myproject.layer3_out_1262_U.if_write & AESL_inst_myproject.layer3_out_1262_U.if_full_n;
    assign fifo_intf_2615.fifo_rd_block = 0;
    assign fifo_intf_2615.fifo_wr_block = 0;
    assign fifo_intf_2615.finish = finish;
    csv_file_dump fifo_csv_dumper_2615;
    csv_file_dump cstatus_csv_dumper_2615;
    df_fifo_monitor fifo_monitor_2615;
    df_fifo_intf fifo_intf_2616(clock,reset);
    assign fifo_intf_2616.rd_en = AESL_inst_myproject.layer3_out_1263_U.if_read & AESL_inst_myproject.layer3_out_1263_U.if_empty_n;
    assign fifo_intf_2616.wr_en = AESL_inst_myproject.layer3_out_1263_U.if_write & AESL_inst_myproject.layer3_out_1263_U.if_full_n;
    assign fifo_intf_2616.fifo_rd_block = 0;
    assign fifo_intf_2616.fifo_wr_block = 0;
    assign fifo_intf_2616.finish = finish;
    csv_file_dump fifo_csv_dumper_2616;
    csv_file_dump cstatus_csv_dumper_2616;
    df_fifo_monitor fifo_monitor_2616;
    df_fifo_intf fifo_intf_2617(clock,reset);
    assign fifo_intf_2617.rd_en = AESL_inst_myproject.layer3_out_1264_U.if_read & AESL_inst_myproject.layer3_out_1264_U.if_empty_n;
    assign fifo_intf_2617.wr_en = AESL_inst_myproject.layer3_out_1264_U.if_write & AESL_inst_myproject.layer3_out_1264_U.if_full_n;
    assign fifo_intf_2617.fifo_rd_block = 0;
    assign fifo_intf_2617.fifo_wr_block = 0;
    assign fifo_intf_2617.finish = finish;
    csv_file_dump fifo_csv_dumper_2617;
    csv_file_dump cstatus_csv_dumper_2617;
    df_fifo_monitor fifo_monitor_2617;
    df_fifo_intf fifo_intf_2618(clock,reset);
    assign fifo_intf_2618.rd_en = AESL_inst_myproject.layer3_out_1265_U.if_read & AESL_inst_myproject.layer3_out_1265_U.if_empty_n;
    assign fifo_intf_2618.wr_en = AESL_inst_myproject.layer3_out_1265_U.if_write & AESL_inst_myproject.layer3_out_1265_U.if_full_n;
    assign fifo_intf_2618.fifo_rd_block = 0;
    assign fifo_intf_2618.fifo_wr_block = 0;
    assign fifo_intf_2618.finish = finish;
    csv_file_dump fifo_csv_dumper_2618;
    csv_file_dump cstatus_csv_dumper_2618;
    df_fifo_monitor fifo_monitor_2618;
    df_fifo_intf fifo_intf_2619(clock,reset);
    assign fifo_intf_2619.rd_en = AESL_inst_myproject.layer3_out_1266_U.if_read & AESL_inst_myproject.layer3_out_1266_U.if_empty_n;
    assign fifo_intf_2619.wr_en = AESL_inst_myproject.layer3_out_1266_U.if_write & AESL_inst_myproject.layer3_out_1266_U.if_full_n;
    assign fifo_intf_2619.fifo_rd_block = 0;
    assign fifo_intf_2619.fifo_wr_block = 0;
    assign fifo_intf_2619.finish = finish;
    csv_file_dump fifo_csv_dumper_2619;
    csv_file_dump cstatus_csv_dumper_2619;
    df_fifo_monitor fifo_monitor_2619;
    df_fifo_intf fifo_intf_2620(clock,reset);
    assign fifo_intf_2620.rd_en = AESL_inst_myproject.layer3_out_1267_U.if_read & AESL_inst_myproject.layer3_out_1267_U.if_empty_n;
    assign fifo_intf_2620.wr_en = AESL_inst_myproject.layer3_out_1267_U.if_write & AESL_inst_myproject.layer3_out_1267_U.if_full_n;
    assign fifo_intf_2620.fifo_rd_block = 0;
    assign fifo_intf_2620.fifo_wr_block = 0;
    assign fifo_intf_2620.finish = finish;
    csv_file_dump fifo_csv_dumper_2620;
    csv_file_dump cstatus_csv_dumper_2620;
    df_fifo_monitor fifo_monitor_2620;
    df_fifo_intf fifo_intf_2621(clock,reset);
    assign fifo_intf_2621.rd_en = AESL_inst_myproject.layer3_out_1268_U.if_read & AESL_inst_myproject.layer3_out_1268_U.if_empty_n;
    assign fifo_intf_2621.wr_en = AESL_inst_myproject.layer3_out_1268_U.if_write & AESL_inst_myproject.layer3_out_1268_U.if_full_n;
    assign fifo_intf_2621.fifo_rd_block = 0;
    assign fifo_intf_2621.fifo_wr_block = 0;
    assign fifo_intf_2621.finish = finish;
    csv_file_dump fifo_csv_dumper_2621;
    csv_file_dump cstatus_csv_dumper_2621;
    df_fifo_monitor fifo_monitor_2621;
    df_fifo_intf fifo_intf_2622(clock,reset);
    assign fifo_intf_2622.rd_en = AESL_inst_myproject.layer3_out_1269_U.if_read & AESL_inst_myproject.layer3_out_1269_U.if_empty_n;
    assign fifo_intf_2622.wr_en = AESL_inst_myproject.layer3_out_1269_U.if_write & AESL_inst_myproject.layer3_out_1269_U.if_full_n;
    assign fifo_intf_2622.fifo_rd_block = 0;
    assign fifo_intf_2622.fifo_wr_block = 0;
    assign fifo_intf_2622.finish = finish;
    csv_file_dump fifo_csv_dumper_2622;
    csv_file_dump cstatus_csv_dumper_2622;
    df_fifo_monitor fifo_monitor_2622;
    df_fifo_intf fifo_intf_2623(clock,reset);
    assign fifo_intf_2623.rd_en = AESL_inst_myproject.layer3_out_1270_U.if_read & AESL_inst_myproject.layer3_out_1270_U.if_empty_n;
    assign fifo_intf_2623.wr_en = AESL_inst_myproject.layer3_out_1270_U.if_write & AESL_inst_myproject.layer3_out_1270_U.if_full_n;
    assign fifo_intf_2623.fifo_rd_block = 0;
    assign fifo_intf_2623.fifo_wr_block = 0;
    assign fifo_intf_2623.finish = finish;
    csv_file_dump fifo_csv_dumper_2623;
    csv_file_dump cstatus_csv_dumper_2623;
    df_fifo_monitor fifo_monitor_2623;
    df_fifo_intf fifo_intf_2624(clock,reset);
    assign fifo_intf_2624.rd_en = AESL_inst_myproject.layer3_out_1271_U.if_read & AESL_inst_myproject.layer3_out_1271_U.if_empty_n;
    assign fifo_intf_2624.wr_en = AESL_inst_myproject.layer3_out_1271_U.if_write & AESL_inst_myproject.layer3_out_1271_U.if_full_n;
    assign fifo_intf_2624.fifo_rd_block = 0;
    assign fifo_intf_2624.fifo_wr_block = 0;
    assign fifo_intf_2624.finish = finish;
    csv_file_dump fifo_csv_dumper_2624;
    csv_file_dump cstatus_csv_dumper_2624;
    df_fifo_monitor fifo_monitor_2624;
    df_fifo_intf fifo_intf_2625(clock,reset);
    assign fifo_intf_2625.rd_en = AESL_inst_myproject.layer3_out_1272_U.if_read & AESL_inst_myproject.layer3_out_1272_U.if_empty_n;
    assign fifo_intf_2625.wr_en = AESL_inst_myproject.layer3_out_1272_U.if_write & AESL_inst_myproject.layer3_out_1272_U.if_full_n;
    assign fifo_intf_2625.fifo_rd_block = 0;
    assign fifo_intf_2625.fifo_wr_block = 0;
    assign fifo_intf_2625.finish = finish;
    csv_file_dump fifo_csv_dumper_2625;
    csv_file_dump cstatus_csv_dumper_2625;
    df_fifo_monitor fifo_monitor_2625;
    df_fifo_intf fifo_intf_2626(clock,reset);
    assign fifo_intf_2626.rd_en = AESL_inst_myproject.layer3_out_1273_U.if_read & AESL_inst_myproject.layer3_out_1273_U.if_empty_n;
    assign fifo_intf_2626.wr_en = AESL_inst_myproject.layer3_out_1273_U.if_write & AESL_inst_myproject.layer3_out_1273_U.if_full_n;
    assign fifo_intf_2626.fifo_rd_block = 0;
    assign fifo_intf_2626.fifo_wr_block = 0;
    assign fifo_intf_2626.finish = finish;
    csv_file_dump fifo_csv_dumper_2626;
    csv_file_dump cstatus_csv_dumper_2626;
    df_fifo_monitor fifo_monitor_2626;
    df_fifo_intf fifo_intf_2627(clock,reset);
    assign fifo_intf_2627.rd_en = AESL_inst_myproject.layer3_out_1274_U.if_read & AESL_inst_myproject.layer3_out_1274_U.if_empty_n;
    assign fifo_intf_2627.wr_en = AESL_inst_myproject.layer3_out_1274_U.if_write & AESL_inst_myproject.layer3_out_1274_U.if_full_n;
    assign fifo_intf_2627.fifo_rd_block = 0;
    assign fifo_intf_2627.fifo_wr_block = 0;
    assign fifo_intf_2627.finish = finish;
    csv_file_dump fifo_csv_dumper_2627;
    csv_file_dump cstatus_csv_dumper_2627;
    df_fifo_monitor fifo_monitor_2627;
    df_fifo_intf fifo_intf_2628(clock,reset);
    assign fifo_intf_2628.rd_en = AESL_inst_myproject.layer3_out_1275_U.if_read & AESL_inst_myproject.layer3_out_1275_U.if_empty_n;
    assign fifo_intf_2628.wr_en = AESL_inst_myproject.layer3_out_1275_U.if_write & AESL_inst_myproject.layer3_out_1275_U.if_full_n;
    assign fifo_intf_2628.fifo_rd_block = 0;
    assign fifo_intf_2628.fifo_wr_block = 0;
    assign fifo_intf_2628.finish = finish;
    csv_file_dump fifo_csv_dumper_2628;
    csv_file_dump cstatus_csv_dumper_2628;
    df_fifo_monitor fifo_monitor_2628;
    df_fifo_intf fifo_intf_2629(clock,reset);
    assign fifo_intf_2629.rd_en = AESL_inst_myproject.layer3_out_1276_U.if_read & AESL_inst_myproject.layer3_out_1276_U.if_empty_n;
    assign fifo_intf_2629.wr_en = AESL_inst_myproject.layer3_out_1276_U.if_write & AESL_inst_myproject.layer3_out_1276_U.if_full_n;
    assign fifo_intf_2629.fifo_rd_block = 0;
    assign fifo_intf_2629.fifo_wr_block = 0;
    assign fifo_intf_2629.finish = finish;
    csv_file_dump fifo_csv_dumper_2629;
    csv_file_dump cstatus_csv_dumper_2629;
    df_fifo_monitor fifo_monitor_2629;
    df_fifo_intf fifo_intf_2630(clock,reset);
    assign fifo_intf_2630.rd_en = AESL_inst_myproject.layer3_out_1277_U.if_read & AESL_inst_myproject.layer3_out_1277_U.if_empty_n;
    assign fifo_intf_2630.wr_en = AESL_inst_myproject.layer3_out_1277_U.if_write & AESL_inst_myproject.layer3_out_1277_U.if_full_n;
    assign fifo_intf_2630.fifo_rd_block = 0;
    assign fifo_intf_2630.fifo_wr_block = 0;
    assign fifo_intf_2630.finish = finish;
    csv_file_dump fifo_csv_dumper_2630;
    csv_file_dump cstatus_csv_dumper_2630;
    df_fifo_monitor fifo_monitor_2630;
    df_fifo_intf fifo_intf_2631(clock,reset);
    assign fifo_intf_2631.rd_en = AESL_inst_myproject.layer3_out_1278_U.if_read & AESL_inst_myproject.layer3_out_1278_U.if_empty_n;
    assign fifo_intf_2631.wr_en = AESL_inst_myproject.layer3_out_1278_U.if_write & AESL_inst_myproject.layer3_out_1278_U.if_full_n;
    assign fifo_intf_2631.fifo_rd_block = 0;
    assign fifo_intf_2631.fifo_wr_block = 0;
    assign fifo_intf_2631.finish = finish;
    csv_file_dump fifo_csv_dumper_2631;
    csv_file_dump cstatus_csv_dumper_2631;
    df_fifo_monitor fifo_monitor_2631;
    df_fifo_intf fifo_intf_2632(clock,reset);
    assign fifo_intf_2632.rd_en = AESL_inst_myproject.layer3_out_1279_U.if_read & AESL_inst_myproject.layer3_out_1279_U.if_empty_n;
    assign fifo_intf_2632.wr_en = AESL_inst_myproject.layer3_out_1279_U.if_write & AESL_inst_myproject.layer3_out_1279_U.if_full_n;
    assign fifo_intf_2632.fifo_rd_block = 0;
    assign fifo_intf_2632.fifo_wr_block = 0;
    assign fifo_intf_2632.finish = finish;
    csv_file_dump fifo_csv_dumper_2632;
    csv_file_dump cstatus_csv_dumper_2632;
    df_fifo_monitor fifo_monitor_2632;
    df_fifo_intf fifo_intf_2633(clock,reset);
    assign fifo_intf_2633.rd_en = AESL_inst_myproject.layer3_out_1280_U.if_read & AESL_inst_myproject.layer3_out_1280_U.if_empty_n;
    assign fifo_intf_2633.wr_en = AESL_inst_myproject.layer3_out_1280_U.if_write & AESL_inst_myproject.layer3_out_1280_U.if_full_n;
    assign fifo_intf_2633.fifo_rd_block = 0;
    assign fifo_intf_2633.fifo_wr_block = 0;
    assign fifo_intf_2633.finish = finish;
    csv_file_dump fifo_csv_dumper_2633;
    csv_file_dump cstatus_csv_dumper_2633;
    df_fifo_monitor fifo_monitor_2633;
    df_fifo_intf fifo_intf_2634(clock,reset);
    assign fifo_intf_2634.rd_en = AESL_inst_myproject.layer3_out_1281_U.if_read & AESL_inst_myproject.layer3_out_1281_U.if_empty_n;
    assign fifo_intf_2634.wr_en = AESL_inst_myproject.layer3_out_1281_U.if_write & AESL_inst_myproject.layer3_out_1281_U.if_full_n;
    assign fifo_intf_2634.fifo_rd_block = 0;
    assign fifo_intf_2634.fifo_wr_block = 0;
    assign fifo_intf_2634.finish = finish;
    csv_file_dump fifo_csv_dumper_2634;
    csv_file_dump cstatus_csv_dumper_2634;
    df_fifo_monitor fifo_monitor_2634;
    df_fifo_intf fifo_intf_2635(clock,reset);
    assign fifo_intf_2635.rd_en = AESL_inst_myproject.layer3_out_1282_U.if_read & AESL_inst_myproject.layer3_out_1282_U.if_empty_n;
    assign fifo_intf_2635.wr_en = AESL_inst_myproject.layer3_out_1282_U.if_write & AESL_inst_myproject.layer3_out_1282_U.if_full_n;
    assign fifo_intf_2635.fifo_rd_block = 0;
    assign fifo_intf_2635.fifo_wr_block = 0;
    assign fifo_intf_2635.finish = finish;
    csv_file_dump fifo_csv_dumper_2635;
    csv_file_dump cstatus_csv_dumper_2635;
    df_fifo_monitor fifo_monitor_2635;
    df_fifo_intf fifo_intf_2636(clock,reset);
    assign fifo_intf_2636.rd_en = AESL_inst_myproject.layer3_out_1283_U.if_read & AESL_inst_myproject.layer3_out_1283_U.if_empty_n;
    assign fifo_intf_2636.wr_en = AESL_inst_myproject.layer3_out_1283_U.if_write & AESL_inst_myproject.layer3_out_1283_U.if_full_n;
    assign fifo_intf_2636.fifo_rd_block = 0;
    assign fifo_intf_2636.fifo_wr_block = 0;
    assign fifo_intf_2636.finish = finish;
    csv_file_dump fifo_csv_dumper_2636;
    csv_file_dump cstatus_csv_dumper_2636;
    df_fifo_monitor fifo_monitor_2636;
    df_fifo_intf fifo_intf_2637(clock,reset);
    assign fifo_intf_2637.rd_en = AESL_inst_myproject.layer3_out_1284_U.if_read & AESL_inst_myproject.layer3_out_1284_U.if_empty_n;
    assign fifo_intf_2637.wr_en = AESL_inst_myproject.layer3_out_1284_U.if_write & AESL_inst_myproject.layer3_out_1284_U.if_full_n;
    assign fifo_intf_2637.fifo_rd_block = 0;
    assign fifo_intf_2637.fifo_wr_block = 0;
    assign fifo_intf_2637.finish = finish;
    csv_file_dump fifo_csv_dumper_2637;
    csv_file_dump cstatus_csv_dumper_2637;
    df_fifo_monitor fifo_monitor_2637;
    df_fifo_intf fifo_intf_2638(clock,reset);
    assign fifo_intf_2638.rd_en = AESL_inst_myproject.layer3_out_1285_U.if_read & AESL_inst_myproject.layer3_out_1285_U.if_empty_n;
    assign fifo_intf_2638.wr_en = AESL_inst_myproject.layer3_out_1285_U.if_write & AESL_inst_myproject.layer3_out_1285_U.if_full_n;
    assign fifo_intf_2638.fifo_rd_block = 0;
    assign fifo_intf_2638.fifo_wr_block = 0;
    assign fifo_intf_2638.finish = finish;
    csv_file_dump fifo_csv_dumper_2638;
    csv_file_dump cstatus_csv_dumper_2638;
    df_fifo_monitor fifo_monitor_2638;
    df_fifo_intf fifo_intf_2639(clock,reset);
    assign fifo_intf_2639.rd_en = AESL_inst_myproject.layer3_out_1286_U.if_read & AESL_inst_myproject.layer3_out_1286_U.if_empty_n;
    assign fifo_intf_2639.wr_en = AESL_inst_myproject.layer3_out_1286_U.if_write & AESL_inst_myproject.layer3_out_1286_U.if_full_n;
    assign fifo_intf_2639.fifo_rd_block = 0;
    assign fifo_intf_2639.fifo_wr_block = 0;
    assign fifo_intf_2639.finish = finish;
    csv_file_dump fifo_csv_dumper_2639;
    csv_file_dump cstatus_csv_dumper_2639;
    df_fifo_monitor fifo_monitor_2639;
    df_fifo_intf fifo_intf_2640(clock,reset);
    assign fifo_intf_2640.rd_en = AESL_inst_myproject.layer3_out_1287_U.if_read & AESL_inst_myproject.layer3_out_1287_U.if_empty_n;
    assign fifo_intf_2640.wr_en = AESL_inst_myproject.layer3_out_1287_U.if_write & AESL_inst_myproject.layer3_out_1287_U.if_full_n;
    assign fifo_intf_2640.fifo_rd_block = 0;
    assign fifo_intf_2640.fifo_wr_block = 0;
    assign fifo_intf_2640.finish = finish;
    csv_file_dump fifo_csv_dumper_2640;
    csv_file_dump cstatus_csv_dumper_2640;
    df_fifo_monitor fifo_monitor_2640;
    df_fifo_intf fifo_intf_2641(clock,reset);
    assign fifo_intf_2641.rd_en = AESL_inst_myproject.layer3_out_1288_U.if_read & AESL_inst_myproject.layer3_out_1288_U.if_empty_n;
    assign fifo_intf_2641.wr_en = AESL_inst_myproject.layer3_out_1288_U.if_write & AESL_inst_myproject.layer3_out_1288_U.if_full_n;
    assign fifo_intf_2641.fifo_rd_block = 0;
    assign fifo_intf_2641.fifo_wr_block = 0;
    assign fifo_intf_2641.finish = finish;
    csv_file_dump fifo_csv_dumper_2641;
    csv_file_dump cstatus_csv_dumper_2641;
    df_fifo_monitor fifo_monitor_2641;
    df_fifo_intf fifo_intf_2642(clock,reset);
    assign fifo_intf_2642.rd_en = AESL_inst_myproject.layer3_out_1289_U.if_read & AESL_inst_myproject.layer3_out_1289_U.if_empty_n;
    assign fifo_intf_2642.wr_en = AESL_inst_myproject.layer3_out_1289_U.if_write & AESL_inst_myproject.layer3_out_1289_U.if_full_n;
    assign fifo_intf_2642.fifo_rd_block = 0;
    assign fifo_intf_2642.fifo_wr_block = 0;
    assign fifo_intf_2642.finish = finish;
    csv_file_dump fifo_csv_dumper_2642;
    csv_file_dump cstatus_csv_dumper_2642;
    df_fifo_monitor fifo_monitor_2642;
    df_fifo_intf fifo_intf_2643(clock,reset);
    assign fifo_intf_2643.rd_en = AESL_inst_myproject.layer3_out_1290_U.if_read & AESL_inst_myproject.layer3_out_1290_U.if_empty_n;
    assign fifo_intf_2643.wr_en = AESL_inst_myproject.layer3_out_1290_U.if_write & AESL_inst_myproject.layer3_out_1290_U.if_full_n;
    assign fifo_intf_2643.fifo_rd_block = 0;
    assign fifo_intf_2643.fifo_wr_block = 0;
    assign fifo_intf_2643.finish = finish;
    csv_file_dump fifo_csv_dumper_2643;
    csv_file_dump cstatus_csv_dumper_2643;
    df_fifo_monitor fifo_monitor_2643;
    df_fifo_intf fifo_intf_2644(clock,reset);
    assign fifo_intf_2644.rd_en = AESL_inst_myproject.layer3_out_1291_U.if_read & AESL_inst_myproject.layer3_out_1291_U.if_empty_n;
    assign fifo_intf_2644.wr_en = AESL_inst_myproject.layer3_out_1291_U.if_write & AESL_inst_myproject.layer3_out_1291_U.if_full_n;
    assign fifo_intf_2644.fifo_rd_block = 0;
    assign fifo_intf_2644.fifo_wr_block = 0;
    assign fifo_intf_2644.finish = finish;
    csv_file_dump fifo_csv_dumper_2644;
    csv_file_dump cstatus_csv_dumper_2644;
    df_fifo_monitor fifo_monitor_2644;
    df_fifo_intf fifo_intf_2645(clock,reset);
    assign fifo_intf_2645.rd_en = AESL_inst_myproject.layer3_out_1292_U.if_read & AESL_inst_myproject.layer3_out_1292_U.if_empty_n;
    assign fifo_intf_2645.wr_en = AESL_inst_myproject.layer3_out_1292_U.if_write & AESL_inst_myproject.layer3_out_1292_U.if_full_n;
    assign fifo_intf_2645.fifo_rd_block = 0;
    assign fifo_intf_2645.fifo_wr_block = 0;
    assign fifo_intf_2645.finish = finish;
    csv_file_dump fifo_csv_dumper_2645;
    csv_file_dump cstatus_csv_dumper_2645;
    df_fifo_monitor fifo_monitor_2645;
    df_fifo_intf fifo_intf_2646(clock,reset);
    assign fifo_intf_2646.rd_en = AESL_inst_myproject.layer3_out_1293_U.if_read & AESL_inst_myproject.layer3_out_1293_U.if_empty_n;
    assign fifo_intf_2646.wr_en = AESL_inst_myproject.layer3_out_1293_U.if_write & AESL_inst_myproject.layer3_out_1293_U.if_full_n;
    assign fifo_intf_2646.fifo_rd_block = 0;
    assign fifo_intf_2646.fifo_wr_block = 0;
    assign fifo_intf_2646.finish = finish;
    csv_file_dump fifo_csv_dumper_2646;
    csv_file_dump cstatus_csv_dumper_2646;
    df_fifo_monitor fifo_monitor_2646;
    df_fifo_intf fifo_intf_2647(clock,reset);
    assign fifo_intf_2647.rd_en = AESL_inst_myproject.layer3_out_1294_U.if_read & AESL_inst_myproject.layer3_out_1294_U.if_empty_n;
    assign fifo_intf_2647.wr_en = AESL_inst_myproject.layer3_out_1294_U.if_write & AESL_inst_myproject.layer3_out_1294_U.if_full_n;
    assign fifo_intf_2647.fifo_rd_block = 0;
    assign fifo_intf_2647.fifo_wr_block = 0;
    assign fifo_intf_2647.finish = finish;
    csv_file_dump fifo_csv_dumper_2647;
    csv_file_dump cstatus_csv_dumper_2647;
    df_fifo_monitor fifo_monitor_2647;
    df_fifo_intf fifo_intf_2648(clock,reset);
    assign fifo_intf_2648.rd_en = AESL_inst_myproject.layer3_out_1295_U.if_read & AESL_inst_myproject.layer3_out_1295_U.if_empty_n;
    assign fifo_intf_2648.wr_en = AESL_inst_myproject.layer3_out_1295_U.if_write & AESL_inst_myproject.layer3_out_1295_U.if_full_n;
    assign fifo_intf_2648.fifo_rd_block = 0;
    assign fifo_intf_2648.fifo_wr_block = 0;
    assign fifo_intf_2648.finish = finish;
    csv_file_dump fifo_csv_dumper_2648;
    csv_file_dump cstatus_csv_dumper_2648;
    df_fifo_monitor fifo_monitor_2648;
    df_fifo_intf fifo_intf_2649(clock,reset);
    assign fifo_intf_2649.rd_en = AESL_inst_myproject.layer3_out_1296_U.if_read & AESL_inst_myproject.layer3_out_1296_U.if_empty_n;
    assign fifo_intf_2649.wr_en = AESL_inst_myproject.layer3_out_1296_U.if_write & AESL_inst_myproject.layer3_out_1296_U.if_full_n;
    assign fifo_intf_2649.fifo_rd_block = 0;
    assign fifo_intf_2649.fifo_wr_block = 0;
    assign fifo_intf_2649.finish = finish;
    csv_file_dump fifo_csv_dumper_2649;
    csv_file_dump cstatus_csv_dumper_2649;
    df_fifo_monitor fifo_monitor_2649;
    df_fifo_intf fifo_intf_2650(clock,reset);
    assign fifo_intf_2650.rd_en = AESL_inst_myproject.layer3_out_1297_U.if_read & AESL_inst_myproject.layer3_out_1297_U.if_empty_n;
    assign fifo_intf_2650.wr_en = AESL_inst_myproject.layer3_out_1297_U.if_write & AESL_inst_myproject.layer3_out_1297_U.if_full_n;
    assign fifo_intf_2650.fifo_rd_block = 0;
    assign fifo_intf_2650.fifo_wr_block = 0;
    assign fifo_intf_2650.finish = finish;
    csv_file_dump fifo_csv_dumper_2650;
    csv_file_dump cstatus_csv_dumper_2650;
    df_fifo_monitor fifo_monitor_2650;
    df_fifo_intf fifo_intf_2651(clock,reset);
    assign fifo_intf_2651.rd_en = AESL_inst_myproject.layer3_out_1298_U.if_read & AESL_inst_myproject.layer3_out_1298_U.if_empty_n;
    assign fifo_intf_2651.wr_en = AESL_inst_myproject.layer3_out_1298_U.if_write & AESL_inst_myproject.layer3_out_1298_U.if_full_n;
    assign fifo_intf_2651.fifo_rd_block = 0;
    assign fifo_intf_2651.fifo_wr_block = 0;
    assign fifo_intf_2651.finish = finish;
    csv_file_dump fifo_csv_dumper_2651;
    csv_file_dump cstatus_csv_dumper_2651;
    df_fifo_monitor fifo_monitor_2651;
    df_fifo_intf fifo_intf_2652(clock,reset);
    assign fifo_intf_2652.rd_en = AESL_inst_myproject.layer3_out_1299_U.if_read & AESL_inst_myproject.layer3_out_1299_U.if_empty_n;
    assign fifo_intf_2652.wr_en = AESL_inst_myproject.layer3_out_1299_U.if_write & AESL_inst_myproject.layer3_out_1299_U.if_full_n;
    assign fifo_intf_2652.fifo_rd_block = 0;
    assign fifo_intf_2652.fifo_wr_block = 0;
    assign fifo_intf_2652.finish = finish;
    csv_file_dump fifo_csv_dumper_2652;
    csv_file_dump cstatus_csv_dumper_2652;
    df_fifo_monitor fifo_monitor_2652;
    df_fifo_intf fifo_intf_2653(clock,reset);
    assign fifo_intf_2653.rd_en = AESL_inst_myproject.layer3_out_1300_U.if_read & AESL_inst_myproject.layer3_out_1300_U.if_empty_n;
    assign fifo_intf_2653.wr_en = AESL_inst_myproject.layer3_out_1300_U.if_write & AESL_inst_myproject.layer3_out_1300_U.if_full_n;
    assign fifo_intf_2653.fifo_rd_block = 0;
    assign fifo_intf_2653.fifo_wr_block = 0;
    assign fifo_intf_2653.finish = finish;
    csv_file_dump fifo_csv_dumper_2653;
    csv_file_dump cstatus_csv_dumper_2653;
    df_fifo_monitor fifo_monitor_2653;
    df_fifo_intf fifo_intf_2654(clock,reset);
    assign fifo_intf_2654.rd_en = AESL_inst_myproject.layer3_out_1301_U.if_read & AESL_inst_myproject.layer3_out_1301_U.if_empty_n;
    assign fifo_intf_2654.wr_en = AESL_inst_myproject.layer3_out_1301_U.if_write & AESL_inst_myproject.layer3_out_1301_U.if_full_n;
    assign fifo_intf_2654.fifo_rd_block = 0;
    assign fifo_intf_2654.fifo_wr_block = 0;
    assign fifo_intf_2654.finish = finish;
    csv_file_dump fifo_csv_dumper_2654;
    csv_file_dump cstatus_csv_dumper_2654;
    df_fifo_monitor fifo_monitor_2654;
    df_fifo_intf fifo_intf_2655(clock,reset);
    assign fifo_intf_2655.rd_en = AESL_inst_myproject.layer3_out_1302_U.if_read & AESL_inst_myproject.layer3_out_1302_U.if_empty_n;
    assign fifo_intf_2655.wr_en = AESL_inst_myproject.layer3_out_1302_U.if_write & AESL_inst_myproject.layer3_out_1302_U.if_full_n;
    assign fifo_intf_2655.fifo_rd_block = 0;
    assign fifo_intf_2655.fifo_wr_block = 0;
    assign fifo_intf_2655.finish = finish;
    csv_file_dump fifo_csv_dumper_2655;
    csv_file_dump cstatus_csv_dumper_2655;
    df_fifo_monitor fifo_monitor_2655;
    df_fifo_intf fifo_intf_2656(clock,reset);
    assign fifo_intf_2656.rd_en = AESL_inst_myproject.layer3_out_1303_U.if_read & AESL_inst_myproject.layer3_out_1303_U.if_empty_n;
    assign fifo_intf_2656.wr_en = AESL_inst_myproject.layer3_out_1303_U.if_write & AESL_inst_myproject.layer3_out_1303_U.if_full_n;
    assign fifo_intf_2656.fifo_rd_block = 0;
    assign fifo_intf_2656.fifo_wr_block = 0;
    assign fifo_intf_2656.finish = finish;
    csv_file_dump fifo_csv_dumper_2656;
    csv_file_dump cstatus_csv_dumper_2656;
    df_fifo_monitor fifo_monitor_2656;
    df_fifo_intf fifo_intf_2657(clock,reset);
    assign fifo_intf_2657.rd_en = AESL_inst_myproject.layer3_out_1304_U.if_read & AESL_inst_myproject.layer3_out_1304_U.if_empty_n;
    assign fifo_intf_2657.wr_en = AESL_inst_myproject.layer3_out_1304_U.if_write & AESL_inst_myproject.layer3_out_1304_U.if_full_n;
    assign fifo_intf_2657.fifo_rd_block = 0;
    assign fifo_intf_2657.fifo_wr_block = 0;
    assign fifo_intf_2657.finish = finish;
    csv_file_dump fifo_csv_dumper_2657;
    csv_file_dump cstatus_csv_dumper_2657;
    df_fifo_monitor fifo_monitor_2657;
    df_fifo_intf fifo_intf_2658(clock,reset);
    assign fifo_intf_2658.rd_en = AESL_inst_myproject.layer3_out_1305_U.if_read & AESL_inst_myproject.layer3_out_1305_U.if_empty_n;
    assign fifo_intf_2658.wr_en = AESL_inst_myproject.layer3_out_1305_U.if_write & AESL_inst_myproject.layer3_out_1305_U.if_full_n;
    assign fifo_intf_2658.fifo_rd_block = 0;
    assign fifo_intf_2658.fifo_wr_block = 0;
    assign fifo_intf_2658.finish = finish;
    csv_file_dump fifo_csv_dumper_2658;
    csv_file_dump cstatus_csv_dumper_2658;
    df_fifo_monitor fifo_monitor_2658;
    df_fifo_intf fifo_intf_2659(clock,reset);
    assign fifo_intf_2659.rd_en = AESL_inst_myproject.layer3_out_1306_U.if_read & AESL_inst_myproject.layer3_out_1306_U.if_empty_n;
    assign fifo_intf_2659.wr_en = AESL_inst_myproject.layer3_out_1306_U.if_write & AESL_inst_myproject.layer3_out_1306_U.if_full_n;
    assign fifo_intf_2659.fifo_rd_block = 0;
    assign fifo_intf_2659.fifo_wr_block = 0;
    assign fifo_intf_2659.finish = finish;
    csv_file_dump fifo_csv_dumper_2659;
    csv_file_dump cstatus_csv_dumper_2659;
    df_fifo_monitor fifo_monitor_2659;
    df_fifo_intf fifo_intf_2660(clock,reset);
    assign fifo_intf_2660.rd_en = AESL_inst_myproject.layer3_out_1307_U.if_read & AESL_inst_myproject.layer3_out_1307_U.if_empty_n;
    assign fifo_intf_2660.wr_en = AESL_inst_myproject.layer3_out_1307_U.if_write & AESL_inst_myproject.layer3_out_1307_U.if_full_n;
    assign fifo_intf_2660.fifo_rd_block = 0;
    assign fifo_intf_2660.fifo_wr_block = 0;
    assign fifo_intf_2660.finish = finish;
    csv_file_dump fifo_csv_dumper_2660;
    csv_file_dump cstatus_csv_dumper_2660;
    df_fifo_monitor fifo_monitor_2660;
    df_fifo_intf fifo_intf_2661(clock,reset);
    assign fifo_intf_2661.rd_en = AESL_inst_myproject.layer3_out_1308_U.if_read & AESL_inst_myproject.layer3_out_1308_U.if_empty_n;
    assign fifo_intf_2661.wr_en = AESL_inst_myproject.layer3_out_1308_U.if_write & AESL_inst_myproject.layer3_out_1308_U.if_full_n;
    assign fifo_intf_2661.fifo_rd_block = 0;
    assign fifo_intf_2661.fifo_wr_block = 0;
    assign fifo_intf_2661.finish = finish;
    csv_file_dump fifo_csv_dumper_2661;
    csv_file_dump cstatus_csv_dumper_2661;
    df_fifo_monitor fifo_monitor_2661;
    df_fifo_intf fifo_intf_2662(clock,reset);
    assign fifo_intf_2662.rd_en = AESL_inst_myproject.layer3_out_1309_U.if_read & AESL_inst_myproject.layer3_out_1309_U.if_empty_n;
    assign fifo_intf_2662.wr_en = AESL_inst_myproject.layer3_out_1309_U.if_write & AESL_inst_myproject.layer3_out_1309_U.if_full_n;
    assign fifo_intf_2662.fifo_rd_block = 0;
    assign fifo_intf_2662.fifo_wr_block = 0;
    assign fifo_intf_2662.finish = finish;
    csv_file_dump fifo_csv_dumper_2662;
    csv_file_dump cstatus_csv_dumper_2662;
    df_fifo_monitor fifo_monitor_2662;
    df_fifo_intf fifo_intf_2663(clock,reset);
    assign fifo_intf_2663.rd_en = AESL_inst_myproject.layer3_out_1310_U.if_read & AESL_inst_myproject.layer3_out_1310_U.if_empty_n;
    assign fifo_intf_2663.wr_en = AESL_inst_myproject.layer3_out_1310_U.if_write & AESL_inst_myproject.layer3_out_1310_U.if_full_n;
    assign fifo_intf_2663.fifo_rd_block = 0;
    assign fifo_intf_2663.fifo_wr_block = 0;
    assign fifo_intf_2663.finish = finish;
    csv_file_dump fifo_csv_dumper_2663;
    csv_file_dump cstatus_csv_dumper_2663;
    df_fifo_monitor fifo_monitor_2663;
    df_fifo_intf fifo_intf_2664(clock,reset);
    assign fifo_intf_2664.rd_en = AESL_inst_myproject.layer3_out_1311_U.if_read & AESL_inst_myproject.layer3_out_1311_U.if_empty_n;
    assign fifo_intf_2664.wr_en = AESL_inst_myproject.layer3_out_1311_U.if_write & AESL_inst_myproject.layer3_out_1311_U.if_full_n;
    assign fifo_intf_2664.fifo_rd_block = 0;
    assign fifo_intf_2664.fifo_wr_block = 0;
    assign fifo_intf_2664.finish = finish;
    csv_file_dump fifo_csv_dumper_2664;
    csv_file_dump cstatus_csv_dumper_2664;
    df_fifo_monitor fifo_monitor_2664;
    df_fifo_intf fifo_intf_2665(clock,reset);
    assign fifo_intf_2665.rd_en = AESL_inst_myproject.layer3_out_1312_U.if_read & AESL_inst_myproject.layer3_out_1312_U.if_empty_n;
    assign fifo_intf_2665.wr_en = AESL_inst_myproject.layer3_out_1312_U.if_write & AESL_inst_myproject.layer3_out_1312_U.if_full_n;
    assign fifo_intf_2665.fifo_rd_block = 0;
    assign fifo_intf_2665.fifo_wr_block = 0;
    assign fifo_intf_2665.finish = finish;
    csv_file_dump fifo_csv_dumper_2665;
    csv_file_dump cstatus_csv_dumper_2665;
    df_fifo_monitor fifo_monitor_2665;
    df_fifo_intf fifo_intf_2666(clock,reset);
    assign fifo_intf_2666.rd_en = AESL_inst_myproject.layer3_out_1313_U.if_read & AESL_inst_myproject.layer3_out_1313_U.if_empty_n;
    assign fifo_intf_2666.wr_en = AESL_inst_myproject.layer3_out_1313_U.if_write & AESL_inst_myproject.layer3_out_1313_U.if_full_n;
    assign fifo_intf_2666.fifo_rd_block = 0;
    assign fifo_intf_2666.fifo_wr_block = 0;
    assign fifo_intf_2666.finish = finish;
    csv_file_dump fifo_csv_dumper_2666;
    csv_file_dump cstatus_csv_dumper_2666;
    df_fifo_monitor fifo_monitor_2666;
    df_fifo_intf fifo_intf_2667(clock,reset);
    assign fifo_intf_2667.rd_en = AESL_inst_myproject.layer3_out_1314_U.if_read & AESL_inst_myproject.layer3_out_1314_U.if_empty_n;
    assign fifo_intf_2667.wr_en = AESL_inst_myproject.layer3_out_1314_U.if_write & AESL_inst_myproject.layer3_out_1314_U.if_full_n;
    assign fifo_intf_2667.fifo_rd_block = 0;
    assign fifo_intf_2667.fifo_wr_block = 0;
    assign fifo_intf_2667.finish = finish;
    csv_file_dump fifo_csv_dumper_2667;
    csv_file_dump cstatus_csv_dumper_2667;
    df_fifo_monitor fifo_monitor_2667;
    df_fifo_intf fifo_intf_2668(clock,reset);
    assign fifo_intf_2668.rd_en = AESL_inst_myproject.layer3_out_1315_U.if_read & AESL_inst_myproject.layer3_out_1315_U.if_empty_n;
    assign fifo_intf_2668.wr_en = AESL_inst_myproject.layer3_out_1315_U.if_write & AESL_inst_myproject.layer3_out_1315_U.if_full_n;
    assign fifo_intf_2668.fifo_rd_block = 0;
    assign fifo_intf_2668.fifo_wr_block = 0;
    assign fifo_intf_2668.finish = finish;
    csv_file_dump fifo_csv_dumper_2668;
    csv_file_dump cstatus_csv_dumper_2668;
    df_fifo_monitor fifo_monitor_2668;
    df_fifo_intf fifo_intf_2669(clock,reset);
    assign fifo_intf_2669.rd_en = AESL_inst_myproject.layer3_out_1316_U.if_read & AESL_inst_myproject.layer3_out_1316_U.if_empty_n;
    assign fifo_intf_2669.wr_en = AESL_inst_myproject.layer3_out_1316_U.if_write & AESL_inst_myproject.layer3_out_1316_U.if_full_n;
    assign fifo_intf_2669.fifo_rd_block = 0;
    assign fifo_intf_2669.fifo_wr_block = 0;
    assign fifo_intf_2669.finish = finish;
    csv_file_dump fifo_csv_dumper_2669;
    csv_file_dump cstatus_csv_dumper_2669;
    df_fifo_monitor fifo_monitor_2669;
    df_fifo_intf fifo_intf_2670(clock,reset);
    assign fifo_intf_2670.rd_en = AESL_inst_myproject.layer3_out_1317_U.if_read & AESL_inst_myproject.layer3_out_1317_U.if_empty_n;
    assign fifo_intf_2670.wr_en = AESL_inst_myproject.layer3_out_1317_U.if_write & AESL_inst_myproject.layer3_out_1317_U.if_full_n;
    assign fifo_intf_2670.fifo_rd_block = 0;
    assign fifo_intf_2670.fifo_wr_block = 0;
    assign fifo_intf_2670.finish = finish;
    csv_file_dump fifo_csv_dumper_2670;
    csv_file_dump cstatus_csv_dumper_2670;
    df_fifo_monitor fifo_monitor_2670;
    df_fifo_intf fifo_intf_2671(clock,reset);
    assign fifo_intf_2671.rd_en = AESL_inst_myproject.layer3_out_1318_U.if_read & AESL_inst_myproject.layer3_out_1318_U.if_empty_n;
    assign fifo_intf_2671.wr_en = AESL_inst_myproject.layer3_out_1318_U.if_write & AESL_inst_myproject.layer3_out_1318_U.if_full_n;
    assign fifo_intf_2671.fifo_rd_block = 0;
    assign fifo_intf_2671.fifo_wr_block = 0;
    assign fifo_intf_2671.finish = finish;
    csv_file_dump fifo_csv_dumper_2671;
    csv_file_dump cstatus_csv_dumper_2671;
    df_fifo_monitor fifo_monitor_2671;
    df_fifo_intf fifo_intf_2672(clock,reset);
    assign fifo_intf_2672.rd_en = AESL_inst_myproject.layer3_out_1319_U.if_read & AESL_inst_myproject.layer3_out_1319_U.if_empty_n;
    assign fifo_intf_2672.wr_en = AESL_inst_myproject.layer3_out_1319_U.if_write & AESL_inst_myproject.layer3_out_1319_U.if_full_n;
    assign fifo_intf_2672.fifo_rd_block = 0;
    assign fifo_intf_2672.fifo_wr_block = 0;
    assign fifo_intf_2672.finish = finish;
    csv_file_dump fifo_csv_dumper_2672;
    csv_file_dump cstatus_csv_dumper_2672;
    df_fifo_monitor fifo_monitor_2672;
    df_fifo_intf fifo_intf_2673(clock,reset);
    assign fifo_intf_2673.rd_en = AESL_inst_myproject.layer3_out_1320_U.if_read & AESL_inst_myproject.layer3_out_1320_U.if_empty_n;
    assign fifo_intf_2673.wr_en = AESL_inst_myproject.layer3_out_1320_U.if_write & AESL_inst_myproject.layer3_out_1320_U.if_full_n;
    assign fifo_intf_2673.fifo_rd_block = 0;
    assign fifo_intf_2673.fifo_wr_block = 0;
    assign fifo_intf_2673.finish = finish;
    csv_file_dump fifo_csv_dumper_2673;
    csv_file_dump cstatus_csv_dumper_2673;
    df_fifo_monitor fifo_monitor_2673;
    df_fifo_intf fifo_intf_2674(clock,reset);
    assign fifo_intf_2674.rd_en = AESL_inst_myproject.layer3_out_1321_U.if_read & AESL_inst_myproject.layer3_out_1321_U.if_empty_n;
    assign fifo_intf_2674.wr_en = AESL_inst_myproject.layer3_out_1321_U.if_write & AESL_inst_myproject.layer3_out_1321_U.if_full_n;
    assign fifo_intf_2674.fifo_rd_block = 0;
    assign fifo_intf_2674.fifo_wr_block = 0;
    assign fifo_intf_2674.finish = finish;
    csv_file_dump fifo_csv_dumper_2674;
    csv_file_dump cstatus_csv_dumper_2674;
    df_fifo_monitor fifo_monitor_2674;
    df_fifo_intf fifo_intf_2675(clock,reset);
    assign fifo_intf_2675.rd_en = AESL_inst_myproject.layer3_out_1322_U.if_read & AESL_inst_myproject.layer3_out_1322_U.if_empty_n;
    assign fifo_intf_2675.wr_en = AESL_inst_myproject.layer3_out_1322_U.if_write & AESL_inst_myproject.layer3_out_1322_U.if_full_n;
    assign fifo_intf_2675.fifo_rd_block = 0;
    assign fifo_intf_2675.fifo_wr_block = 0;
    assign fifo_intf_2675.finish = finish;
    csv_file_dump fifo_csv_dumper_2675;
    csv_file_dump cstatus_csv_dumper_2675;
    df_fifo_monitor fifo_monitor_2675;
    df_fifo_intf fifo_intf_2676(clock,reset);
    assign fifo_intf_2676.rd_en = AESL_inst_myproject.layer3_out_1323_U.if_read & AESL_inst_myproject.layer3_out_1323_U.if_empty_n;
    assign fifo_intf_2676.wr_en = AESL_inst_myproject.layer3_out_1323_U.if_write & AESL_inst_myproject.layer3_out_1323_U.if_full_n;
    assign fifo_intf_2676.fifo_rd_block = 0;
    assign fifo_intf_2676.fifo_wr_block = 0;
    assign fifo_intf_2676.finish = finish;
    csv_file_dump fifo_csv_dumper_2676;
    csv_file_dump cstatus_csv_dumper_2676;
    df_fifo_monitor fifo_monitor_2676;
    df_fifo_intf fifo_intf_2677(clock,reset);
    assign fifo_intf_2677.rd_en = AESL_inst_myproject.layer3_out_1324_U.if_read & AESL_inst_myproject.layer3_out_1324_U.if_empty_n;
    assign fifo_intf_2677.wr_en = AESL_inst_myproject.layer3_out_1324_U.if_write & AESL_inst_myproject.layer3_out_1324_U.if_full_n;
    assign fifo_intf_2677.fifo_rd_block = 0;
    assign fifo_intf_2677.fifo_wr_block = 0;
    assign fifo_intf_2677.finish = finish;
    csv_file_dump fifo_csv_dumper_2677;
    csv_file_dump cstatus_csv_dumper_2677;
    df_fifo_monitor fifo_monitor_2677;
    df_fifo_intf fifo_intf_2678(clock,reset);
    assign fifo_intf_2678.rd_en = AESL_inst_myproject.layer3_out_1325_U.if_read & AESL_inst_myproject.layer3_out_1325_U.if_empty_n;
    assign fifo_intf_2678.wr_en = AESL_inst_myproject.layer3_out_1325_U.if_write & AESL_inst_myproject.layer3_out_1325_U.if_full_n;
    assign fifo_intf_2678.fifo_rd_block = 0;
    assign fifo_intf_2678.fifo_wr_block = 0;
    assign fifo_intf_2678.finish = finish;
    csv_file_dump fifo_csv_dumper_2678;
    csv_file_dump cstatus_csv_dumper_2678;
    df_fifo_monitor fifo_monitor_2678;
    df_fifo_intf fifo_intf_2679(clock,reset);
    assign fifo_intf_2679.rd_en = AESL_inst_myproject.layer3_out_1326_U.if_read & AESL_inst_myproject.layer3_out_1326_U.if_empty_n;
    assign fifo_intf_2679.wr_en = AESL_inst_myproject.layer3_out_1326_U.if_write & AESL_inst_myproject.layer3_out_1326_U.if_full_n;
    assign fifo_intf_2679.fifo_rd_block = 0;
    assign fifo_intf_2679.fifo_wr_block = 0;
    assign fifo_intf_2679.finish = finish;
    csv_file_dump fifo_csv_dumper_2679;
    csv_file_dump cstatus_csv_dumper_2679;
    df_fifo_monitor fifo_monitor_2679;
    df_fifo_intf fifo_intf_2680(clock,reset);
    assign fifo_intf_2680.rd_en = AESL_inst_myproject.layer3_out_1327_U.if_read & AESL_inst_myproject.layer3_out_1327_U.if_empty_n;
    assign fifo_intf_2680.wr_en = AESL_inst_myproject.layer3_out_1327_U.if_write & AESL_inst_myproject.layer3_out_1327_U.if_full_n;
    assign fifo_intf_2680.fifo_rd_block = 0;
    assign fifo_intf_2680.fifo_wr_block = 0;
    assign fifo_intf_2680.finish = finish;
    csv_file_dump fifo_csv_dumper_2680;
    csv_file_dump cstatus_csv_dumper_2680;
    df_fifo_monitor fifo_monitor_2680;
    df_fifo_intf fifo_intf_2681(clock,reset);
    assign fifo_intf_2681.rd_en = AESL_inst_myproject.layer3_out_1328_U.if_read & AESL_inst_myproject.layer3_out_1328_U.if_empty_n;
    assign fifo_intf_2681.wr_en = AESL_inst_myproject.layer3_out_1328_U.if_write & AESL_inst_myproject.layer3_out_1328_U.if_full_n;
    assign fifo_intf_2681.fifo_rd_block = 0;
    assign fifo_intf_2681.fifo_wr_block = 0;
    assign fifo_intf_2681.finish = finish;
    csv_file_dump fifo_csv_dumper_2681;
    csv_file_dump cstatus_csv_dumper_2681;
    df_fifo_monitor fifo_monitor_2681;
    df_fifo_intf fifo_intf_2682(clock,reset);
    assign fifo_intf_2682.rd_en = AESL_inst_myproject.layer3_out_1329_U.if_read & AESL_inst_myproject.layer3_out_1329_U.if_empty_n;
    assign fifo_intf_2682.wr_en = AESL_inst_myproject.layer3_out_1329_U.if_write & AESL_inst_myproject.layer3_out_1329_U.if_full_n;
    assign fifo_intf_2682.fifo_rd_block = 0;
    assign fifo_intf_2682.fifo_wr_block = 0;
    assign fifo_intf_2682.finish = finish;
    csv_file_dump fifo_csv_dumper_2682;
    csv_file_dump cstatus_csv_dumper_2682;
    df_fifo_monitor fifo_monitor_2682;
    df_fifo_intf fifo_intf_2683(clock,reset);
    assign fifo_intf_2683.rd_en = AESL_inst_myproject.layer3_out_1330_U.if_read & AESL_inst_myproject.layer3_out_1330_U.if_empty_n;
    assign fifo_intf_2683.wr_en = AESL_inst_myproject.layer3_out_1330_U.if_write & AESL_inst_myproject.layer3_out_1330_U.if_full_n;
    assign fifo_intf_2683.fifo_rd_block = 0;
    assign fifo_intf_2683.fifo_wr_block = 0;
    assign fifo_intf_2683.finish = finish;
    csv_file_dump fifo_csv_dumper_2683;
    csv_file_dump cstatus_csv_dumper_2683;
    df_fifo_monitor fifo_monitor_2683;
    df_fifo_intf fifo_intf_2684(clock,reset);
    assign fifo_intf_2684.rd_en = AESL_inst_myproject.layer3_out_1331_U.if_read & AESL_inst_myproject.layer3_out_1331_U.if_empty_n;
    assign fifo_intf_2684.wr_en = AESL_inst_myproject.layer3_out_1331_U.if_write & AESL_inst_myproject.layer3_out_1331_U.if_full_n;
    assign fifo_intf_2684.fifo_rd_block = 0;
    assign fifo_intf_2684.fifo_wr_block = 0;
    assign fifo_intf_2684.finish = finish;
    csv_file_dump fifo_csv_dumper_2684;
    csv_file_dump cstatus_csv_dumper_2684;
    df_fifo_monitor fifo_monitor_2684;
    df_fifo_intf fifo_intf_2685(clock,reset);
    assign fifo_intf_2685.rd_en = AESL_inst_myproject.layer3_out_1332_U.if_read & AESL_inst_myproject.layer3_out_1332_U.if_empty_n;
    assign fifo_intf_2685.wr_en = AESL_inst_myproject.layer3_out_1332_U.if_write & AESL_inst_myproject.layer3_out_1332_U.if_full_n;
    assign fifo_intf_2685.fifo_rd_block = 0;
    assign fifo_intf_2685.fifo_wr_block = 0;
    assign fifo_intf_2685.finish = finish;
    csv_file_dump fifo_csv_dumper_2685;
    csv_file_dump cstatus_csv_dumper_2685;
    df_fifo_monitor fifo_monitor_2685;
    df_fifo_intf fifo_intf_2686(clock,reset);
    assign fifo_intf_2686.rd_en = AESL_inst_myproject.layer3_out_1333_U.if_read & AESL_inst_myproject.layer3_out_1333_U.if_empty_n;
    assign fifo_intf_2686.wr_en = AESL_inst_myproject.layer3_out_1333_U.if_write & AESL_inst_myproject.layer3_out_1333_U.if_full_n;
    assign fifo_intf_2686.fifo_rd_block = 0;
    assign fifo_intf_2686.fifo_wr_block = 0;
    assign fifo_intf_2686.finish = finish;
    csv_file_dump fifo_csv_dumper_2686;
    csv_file_dump cstatus_csv_dumper_2686;
    df_fifo_monitor fifo_monitor_2686;
    df_fifo_intf fifo_intf_2687(clock,reset);
    assign fifo_intf_2687.rd_en = AESL_inst_myproject.layer3_out_1334_U.if_read & AESL_inst_myproject.layer3_out_1334_U.if_empty_n;
    assign fifo_intf_2687.wr_en = AESL_inst_myproject.layer3_out_1334_U.if_write & AESL_inst_myproject.layer3_out_1334_U.if_full_n;
    assign fifo_intf_2687.fifo_rd_block = 0;
    assign fifo_intf_2687.fifo_wr_block = 0;
    assign fifo_intf_2687.finish = finish;
    csv_file_dump fifo_csv_dumper_2687;
    csv_file_dump cstatus_csv_dumper_2687;
    df_fifo_monitor fifo_monitor_2687;
    df_fifo_intf fifo_intf_2688(clock,reset);
    assign fifo_intf_2688.rd_en = AESL_inst_myproject.layer3_out_1335_U.if_read & AESL_inst_myproject.layer3_out_1335_U.if_empty_n;
    assign fifo_intf_2688.wr_en = AESL_inst_myproject.layer3_out_1335_U.if_write & AESL_inst_myproject.layer3_out_1335_U.if_full_n;
    assign fifo_intf_2688.fifo_rd_block = 0;
    assign fifo_intf_2688.fifo_wr_block = 0;
    assign fifo_intf_2688.finish = finish;
    csv_file_dump fifo_csv_dumper_2688;
    csv_file_dump cstatus_csv_dumper_2688;
    df_fifo_monitor fifo_monitor_2688;
    df_fifo_intf fifo_intf_2689(clock,reset);
    assign fifo_intf_2689.rd_en = AESL_inst_myproject.layer3_out_1336_U.if_read & AESL_inst_myproject.layer3_out_1336_U.if_empty_n;
    assign fifo_intf_2689.wr_en = AESL_inst_myproject.layer3_out_1336_U.if_write & AESL_inst_myproject.layer3_out_1336_U.if_full_n;
    assign fifo_intf_2689.fifo_rd_block = 0;
    assign fifo_intf_2689.fifo_wr_block = 0;
    assign fifo_intf_2689.finish = finish;
    csv_file_dump fifo_csv_dumper_2689;
    csv_file_dump cstatus_csv_dumper_2689;
    df_fifo_monitor fifo_monitor_2689;
    df_fifo_intf fifo_intf_2690(clock,reset);
    assign fifo_intf_2690.rd_en = AESL_inst_myproject.layer3_out_1337_U.if_read & AESL_inst_myproject.layer3_out_1337_U.if_empty_n;
    assign fifo_intf_2690.wr_en = AESL_inst_myproject.layer3_out_1337_U.if_write & AESL_inst_myproject.layer3_out_1337_U.if_full_n;
    assign fifo_intf_2690.fifo_rd_block = 0;
    assign fifo_intf_2690.fifo_wr_block = 0;
    assign fifo_intf_2690.finish = finish;
    csv_file_dump fifo_csv_dumper_2690;
    csv_file_dump cstatus_csv_dumper_2690;
    df_fifo_monitor fifo_monitor_2690;
    df_fifo_intf fifo_intf_2691(clock,reset);
    assign fifo_intf_2691.rd_en = AESL_inst_myproject.layer3_out_1338_U.if_read & AESL_inst_myproject.layer3_out_1338_U.if_empty_n;
    assign fifo_intf_2691.wr_en = AESL_inst_myproject.layer3_out_1338_U.if_write & AESL_inst_myproject.layer3_out_1338_U.if_full_n;
    assign fifo_intf_2691.fifo_rd_block = 0;
    assign fifo_intf_2691.fifo_wr_block = 0;
    assign fifo_intf_2691.finish = finish;
    csv_file_dump fifo_csv_dumper_2691;
    csv_file_dump cstatus_csv_dumper_2691;
    df_fifo_monitor fifo_monitor_2691;
    df_fifo_intf fifo_intf_2692(clock,reset);
    assign fifo_intf_2692.rd_en = AESL_inst_myproject.layer3_out_1339_U.if_read & AESL_inst_myproject.layer3_out_1339_U.if_empty_n;
    assign fifo_intf_2692.wr_en = AESL_inst_myproject.layer3_out_1339_U.if_write & AESL_inst_myproject.layer3_out_1339_U.if_full_n;
    assign fifo_intf_2692.fifo_rd_block = 0;
    assign fifo_intf_2692.fifo_wr_block = 0;
    assign fifo_intf_2692.finish = finish;
    csv_file_dump fifo_csv_dumper_2692;
    csv_file_dump cstatus_csv_dumper_2692;
    df_fifo_monitor fifo_monitor_2692;
    df_fifo_intf fifo_intf_2693(clock,reset);
    assign fifo_intf_2693.rd_en = AESL_inst_myproject.layer3_out_1340_U.if_read & AESL_inst_myproject.layer3_out_1340_U.if_empty_n;
    assign fifo_intf_2693.wr_en = AESL_inst_myproject.layer3_out_1340_U.if_write & AESL_inst_myproject.layer3_out_1340_U.if_full_n;
    assign fifo_intf_2693.fifo_rd_block = 0;
    assign fifo_intf_2693.fifo_wr_block = 0;
    assign fifo_intf_2693.finish = finish;
    csv_file_dump fifo_csv_dumper_2693;
    csv_file_dump cstatus_csv_dumper_2693;
    df_fifo_monitor fifo_monitor_2693;
    df_fifo_intf fifo_intf_2694(clock,reset);
    assign fifo_intf_2694.rd_en = AESL_inst_myproject.layer3_out_1341_U.if_read & AESL_inst_myproject.layer3_out_1341_U.if_empty_n;
    assign fifo_intf_2694.wr_en = AESL_inst_myproject.layer3_out_1341_U.if_write & AESL_inst_myproject.layer3_out_1341_U.if_full_n;
    assign fifo_intf_2694.fifo_rd_block = 0;
    assign fifo_intf_2694.fifo_wr_block = 0;
    assign fifo_intf_2694.finish = finish;
    csv_file_dump fifo_csv_dumper_2694;
    csv_file_dump cstatus_csv_dumper_2694;
    df_fifo_monitor fifo_monitor_2694;
    df_fifo_intf fifo_intf_2695(clock,reset);
    assign fifo_intf_2695.rd_en = AESL_inst_myproject.layer3_out_1342_U.if_read & AESL_inst_myproject.layer3_out_1342_U.if_empty_n;
    assign fifo_intf_2695.wr_en = AESL_inst_myproject.layer3_out_1342_U.if_write & AESL_inst_myproject.layer3_out_1342_U.if_full_n;
    assign fifo_intf_2695.fifo_rd_block = 0;
    assign fifo_intf_2695.fifo_wr_block = 0;
    assign fifo_intf_2695.finish = finish;
    csv_file_dump fifo_csv_dumper_2695;
    csv_file_dump cstatus_csv_dumper_2695;
    df_fifo_monitor fifo_monitor_2695;
    df_fifo_intf fifo_intf_2696(clock,reset);
    assign fifo_intf_2696.rd_en = AESL_inst_myproject.layer3_out_1343_U.if_read & AESL_inst_myproject.layer3_out_1343_U.if_empty_n;
    assign fifo_intf_2696.wr_en = AESL_inst_myproject.layer3_out_1343_U.if_write & AESL_inst_myproject.layer3_out_1343_U.if_full_n;
    assign fifo_intf_2696.fifo_rd_block = 0;
    assign fifo_intf_2696.fifo_wr_block = 0;
    assign fifo_intf_2696.finish = finish;
    csv_file_dump fifo_csv_dumper_2696;
    csv_file_dump cstatus_csv_dumper_2696;
    df_fifo_monitor fifo_monitor_2696;
    df_fifo_intf fifo_intf_2697(clock,reset);
    assign fifo_intf_2697.rd_en = AESL_inst_myproject.layer3_out_1344_U.if_read & AESL_inst_myproject.layer3_out_1344_U.if_empty_n;
    assign fifo_intf_2697.wr_en = AESL_inst_myproject.layer3_out_1344_U.if_write & AESL_inst_myproject.layer3_out_1344_U.if_full_n;
    assign fifo_intf_2697.fifo_rd_block = 0;
    assign fifo_intf_2697.fifo_wr_block = 0;
    assign fifo_intf_2697.finish = finish;
    csv_file_dump fifo_csv_dumper_2697;
    csv_file_dump cstatus_csv_dumper_2697;
    df_fifo_monitor fifo_monitor_2697;
    df_fifo_intf fifo_intf_2698(clock,reset);
    assign fifo_intf_2698.rd_en = AESL_inst_myproject.layer3_out_1345_U.if_read & AESL_inst_myproject.layer3_out_1345_U.if_empty_n;
    assign fifo_intf_2698.wr_en = AESL_inst_myproject.layer3_out_1345_U.if_write & AESL_inst_myproject.layer3_out_1345_U.if_full_n;
    assign fifo_intf_2698.fifo_rd_block = 0;
    assign fifo_intf_2698.fifo_wr_block = 0;
    assign fifo_intf_2698.finish = finish;
    csv_file_dump fifo_csv_dumper_2698;
    csv_file_dump cstatus_csv_dumper_2698;
    df_fifo_monitor fifo_monitor_2698;
    df_fifo_intf fifo_intf_2699(clock,reset);
    assign fifo_intf_2699.rd_en = AESL_inst_myproject.layer3_out_1346_U.if_read & AESL_inst_myproject.layer3_out_1346_U.if_empty_n;
    assign fifo_intf_2699.wr_en = AESL_inst_myproject.layer3_out_1346_U.if_write & AESL_inst_myproject.layer3_out_1346_U.if_full_n;
    assign fifo_intf_2699.fifo_rd_block = 0;
    assign fifo_intf_2699.fifo_wr_block = 0;
    assign fifo_intf_2699.finish = finish;
    csv_file_dump fifo_csv_dumper_2699;
    csv_file_dump cstatus_csv_dumper_2699;
    df_fifo_monitor fifo_monitor_2699;
    df_fifo_intf fifo_intf_2700(clock,reset);
    assign fifo_intf_2700.rd_en = AESL_inst_myproject.layer3_out_1347_U.if_read & AESL_inst_myproject.layer3_out_1347_U.if_empty_n;
    assign fifo_intf_2700.wr_en = AESL_inst_myproject.layer3_out_1347_U.if_write & AESL_inst_myproject.layer3_out_1347_U.if_full_n;
    assign fifo_intf_2700.fifo_rd_block = 0;
    assign fifo_intf_2700.fifo_wr_block = 0;
    assign fifo_intf_2700.finish = finish;
    csv_file_dump fifo_csv_dumper_2700;
    csv_file_dump cstatus_csv_dumper_2700;
    df_fifo_monitor fifo_monitor_2700;
    df_fifo_intf fifo_intf_2701(clock,reset);
    assign fifo_intf_2701.rd_en = AESL_inst_myproject.layer3_out_1348_U.if_read & AESL_inst_myproject.layer3_out_1348_U.if_empty_n;
    assign fifo_intf_2701.wr_en = AESL_inst_myproject.layer3_out_1348_U.if_write & AESL_inst_myproject.layer3_out_1348_U.if_full_n;
    assign fifo_intf_2701.fifo_rd_block = 0;
    assign fifo_intf_2701.fifo_wr_block = 0;
    assign fifo_intf_2701.finish = finish;
    csv_file_dump fifo_csv_dumper_2701;
    csv_file_dump cstatus_csv_dumper_2701;
    df_fifo_monitor fifo_monitor_2701;
    df_fifo_intf fifo_intf_2702(clock,reset);
    assign fifo_intf_2702.rd_en = AESL_inst_myproject.layer3_out_1349_U.if_read & AESL_inst_myproject.layer3_out_1349_U.if_empty_n;
    assign fifo_intf_2702.wr_en = AESL_inst_myproject.layer3_out_1349_U.if_write & AESL_inst_myproject.layer3_out_1349_U.if_full_n;
    assign fifo_intf_2702.fifo_rd_block = 0;
    assign fifo_intf_2702.fifo_wr_block = 0;
    assign fifo_intf_2702.finish = finish;
    csv_file_dump fifo_csv_dumper_2702;
    csv_file_dump cstatus_csv_dumper_2702;
    df_fifo_monitor fifo_monitor_2702;
    df_fifo_intf fifo_intf_2703(clock,reset);
    assign fifo_intf_2703.rd_en = AESL_inst_myproject.layer3_out_1350_U.if_read & AESL_inst_myproject.layer3_out_1350_U.if_empty_n;
    assign fifo_intf_2703.wr_en = AESL_inst_myproject.layer3_out_1350_U.if_write & AESL_inst_myproject.layer3_out_1350_U.if_full_n;
    assign fifo_intf_2703.fifo_rd_block = 0;
    assign fifo_intf_2703.fifo_wr_block = 0;
    assign fifo_intf_2703.finish = finish;
    csv_file_dump fifo_csv_dumper_2703;
    csv_file_dump cstatus_csv_dumper_2703;
    df_fifo_monitor fifo_monitor_2703;
    df_fifo_intf fifo_intf_2704(clock,reset);
    assign fifo_intf_2704.rd_en = AESL_inst_myproject.layer3_out_1351_U.if_read & AESL_inst_myproject.layer3_out_1351_U.if_empty_n;
    assign fifo_intf_2704.wr_en = AESL_inst_myproject.layer3_out_1351_U.if_write & AESL_inst_myproject.layer3_out_1351_U.if_full_n;
    assign fifo_intf_2704.fifo_rd_block = 0;
    assign fifo_intf_2704.fifo_wr_block = 0;
    assign fifo_intf_2704.finish = finish;
    csv_file_dump fifo_csv_dumper_2704;
    csv_file_dump cstatus_csv_dumper_2704;
    df_fifo_monitor fifo_monitor_2704;
    df_fifo_intf fifo_intf_2705(clock,reset);
    assign fifo_intf_2705.rd_en = AESL_inst_myproject.layer5_out_U.if_read & AESL_inst_myproject.layer5_out_U.if_empty_n;
    assign fifo_intf_2705.wr_en = AESL_inst_myproject.layer5_out_U.if_write & AESL_inst_myproject.layer5_out_U.if_full_n;
    assign fifo_intf_2705.fifo_rd_block = 0;
    assign fifo_intf_2705.fifo_wr_block = 0;
    assign fifo_intf_2705.finish = finish;
    csv_file_dump fifo_csv_dumper_2705;
    csv_file_dump cstatus_csv_dumper_2705;
    df_fifo_monitor fifo_monitor_2705;
    df_fifo_intf fifo_intf_2706(clock,reset);
    assign fifo_intf_2706.rd_en = AESL_inst_myproject.layer5_out_1_U.if_read & AESL_inst_myproject.layer5_out_1_U.if_empty_n;
    assign fifo_intf_2706.wr_en = AESL_inst_myproject.layer5_out_1_U.if_write & AESL_inst_myproject.layer5_out_1_U.if_full_n;
    assign fifo_intf_2706.fifo_rd_block = 0;
    assign fifo_intf_2706.fifo_wr_block = 0;
    assign fifo_intf_2706.finish = finish;
    csv_file_dump fifo_csv_dumper_2706;
    csv_file_dump cstatus_csv_dumper_2706;
    df_fifo_monitor fifo_monitor_2706;
    df_fifo_intf fifo_intf_2707(clock,reset);
    assign fifo_intf_2707.rd_en = AESL_inst_myproject.layer5_out_2_U.if_read & AESL_inst_myproject.layer5_out_2_U.if_empty_n;
    assign fifo_intf_2707.wr_en = AESL_inst_myproject.layer5_out_2_U.if_write & AESL_inst_myproject.layer5_out_2_U.if_full_n;
    assign fifo_intf_2707.fifo_rd_block = 0;
    assign fifo_intf_2707.fifo_wr_block = 0;
    assign fifo_intf_2707.finish = finish;
    csv_file_dump fifo_csv_dumper_2707;
    csv_file_dump cstatus_csv_dumper_2707;
    df_fifo_monitor fifo_monitor_2707;
    df_fifo_intf fifo_intf_2708(clock,reset);
    assign fifo_intf_2708.rd_en = AESL_inst_myproject.layer5_out_3_U.if_read & AESL_inst_myproject.layer5_out_3_U.if_empty_n;
    assign fifo_intf_2708.wr_en = AESL_inst_myproject.layer5_out_3_U.if_write & AESL_inst_myproject.layer5_out_3_U.if_full_n;
    assign fifo_intf_2708.fifo_rd_block = 0;
    assign fifo_intf_2708.fifo_wr_block = 0;
    assign fifo_intf_2708.finish = finish;
    csv_file_dump fifo_csv_dumper_2708;
    csv_file_dump cstatus_csv_dumper_2708;
    df_fifo_monitor fifo_monitor_2708;
    df_fifo_intf fifo_intf_2709(clock,reset);
    assign fifo_intf_2709.rd_en = AESL_inst_myproject.layer5_out_4_U.if_read & AESL_inst_myproject.layer5_out_4_U.if_empty_n;
    assign fifo_intf_2709.wr_en = AESL_inst_myproject.layer5_out_4_U.if_write & AESL_inst_myproject.layer5_out_4_U.if_full_n;
    assign fifo_intf_2709.fifo_rd_block = 0;
    assign fifo_intf_2709.fifo_wr_block = 0;
    assign fifo_intf_2709.finish = finish;
    csv_file_dump fifo_csv_dumper_2709;
    csv_file_dump cstatus_csv_dumper_2709;
    df_fifo_monitor fifo_monitor_2709;
    df_fifo_intf fifo_intf_2710(clock,reset);
    assign fifo_intf_2710.rd_en = AESL_inst_myproject.layer5_out_5_U.if_read & AESL_inst_myproject.layer5_out_5_U.if_empty_n;
    assign fifo_intf_2710.wr_en = AESL_inst_myproject.layer5_out_5_U.if_write & AESL_inst_myproject.layer5_out_5_U.if_full_n;
    assign fifo_intf_2710.fifo_rd_block = 0;
    assign fifo_intf_2710.fifo_wr_block = 0;
    assign fifo_intf_2710.finish = finish;
    csv_file_dump fifo_csv_dumper_2710;
    csv_file_dump cstatus_csv_dumper_2710;
    df_fifo_monitor fifo_monitor_2710;
    df_fifo_intf fifo_intf_2711(clock,reset);
    assign fifo_intf_2711.rd_en = AESL_inst_myproject.layer5_out_6_U.if_read & AESL_inst_myproject.layer5_out_6_U.if_empty_n;
    assign fifo_intf_2711.wr_en = AESL_inst_myproject.layer5_out_6_U.if_write & AESL_inst_myproject.layer5_out_6_U.if_full_n;
    assign fifo_intf_2711.fifo_rd_block = 0;
    assign fifo_intf_2711.fifo_wr_block = 0;
    assign fifo_intf_2711.finish = finish;
    csv_file_dump fifo_csv_dumper_2711;
    csv_file_dump cstatus_csv_dumper_2711;
    df_fifo_monitor fifo_monitor_2711;
    df_fifo_intf fifo_intf_2712(clock,reset);
    assign fifo_intf_2712.rd_en = AESL_inst_myproject.layer5_out_7_U.if_read & AESL_inst_myproject.layer5_out_7_U.if_empty_n;
    assign fifo_intf_2712.wr_en = AESL_inst_myproject.layer5_out_7_U.if_write & AESL_inst_myproject.layer5_out_7_U.if_full_n;
    assign fifo_intf_2712.fifo_rd_block = 0;
    assign fifo_intf_2712.fifo_wr_block = 0;
    assign fifo_intf_2712.finish = finish;
    csv_file_dump fifo_csv_dumper_2712;
    csv_file_dump cstatus_csv_dumper_2712;
    df_fifo_monitor fifo_monitor_2712;
    df_fifo_intf fifo_intf_2713(clock,reset);
    assign fifo_intf_2713.rd_en = AESL_inst_myproject.layer5_out_8_U.if_read & AESL_inst_myproject.layer5_out_8_U.if_empty_n;
    assign fifo_intf_2713.wr_en = AESL_inst_myproject.layer5_out_8_U.if_write & AESL_inst_myproject.layer5_out_8_U.if_full_n;
    assign fifo_intf_2713.fifo_rd_block = 0;
    assign fifo_intf_2713.fifo_wr_block = 0;
    assign fifo_intf_2713.finish = finish;
    csv_file_dump fifo_csv_dumper_2713;
    csv_file_dump cstatus_csv_dumper_2713;
    df_fifo_monitor fifo_monitor_2713;
    df_fifo_intf fifo_intf_2714(clock,reset);
    assign fifo_intf_2714.rd_en = AESL_inst_myproject.layer5_out_9_U.if_read & AESL_inst_myproject.layer5_out_9_U.if_empty_n;
    assign fifo_intf_2714.wr_en = AESL_inst_myproject.layer5_out_9_U.if_write & AESL_inst_myproject.layer5_out_9_U.if_full_n;
    assign fifo_intf_2714.fifo_rd_block = 0;
    assign fifo_intf_2714.fifo_wr_block = 0;
    assign fifo_intf_2714.finish = finish;
    csv_file_dump fifo_csv_dumper_2714;
    csv_file_dump cstatus_csv_dumper_2714;
    df_fifo_monitor fifo_monitor_2714;

logic region_0_idle;
logic [31:0] region_0_start_cnt;
logic [31:0] region_0_done_cnt;
assign region_0_idle = (region_0_start_cnt == region_0_done_cnt) && AESL_inst_myproject.ap_start == 1'b0 ;
always @(posedge clock) begin
    if (reset == 1'b1)
        region_0_start_cnt <= 32'h0;
    else if (AESL_inst_myproject.ap_start == 1'b1 && AESL_inst_myproject.ap_ready == 1'b1)
        region_0_start_cnt <= region_0_start_cnt + 32'h1;
    else;
end
always @(posedge clock) begin
    if (reset == 1'b1)
        region_0_done_cnt <= 32'h0;
    else if (AESL_inst_myproject.ap_done == 1'b1)
        region_0_done_cnt <= region_0_done_cnt + 32'h1;
    else;
end


    df_process_intf process_intf_1(clock,reset);
    assign process_intf_1.ap_start = AESL_inst_myproject.conv_2d_cl_ap_fixed_6_2_5_3_0_ap_fixed_6_2_5_3_0_config2_U0.ap_start;
    assign process_intf_1.ap_ready = AESL_inst_myproject.conv_2d_cl_ap_fixed_6_2_5_3_0_ap_fixed_6_2_5_3_0_config2_U0.ap_ready;
    assign process_intf_1.ap_done = AESL_inst_myproject.conv_2d_cl_ap_fixed_6_2_5_3_0_ap_fixed_6_2_5_3_0_config2_U0.ap_done;
    assign process_intf_1.ap_continue = AESL_inst_myproject.conv_2d_cl_ap_fixed_6_2_5_3_0_ap_fixed_6_2_5_3_0_config2_U0.ap_continue;
    assign process_intf_1.real_start = AESL_inst_myproject.conv_2d_cl_ap_fixed_6_2_5_3_0_ap_fixed_6_2_5_3_0_config2_U0.ap_start;
    assign process_intf_1.pin_stall = 1'b0;
    assign process_intf_1.pout_stall = 1'b0;
    assign process_intf_1.cin_stall = 1'b0;
    assign process_intf_1.cout_stall = 1'b0;
    assign process_intf_1.region_idle = region_0_idle;
    assign process_intf_1.finish = finish;
    csv_file_dump pstall_csv_dumper_1;
    csv_file_dump pstatus_csv_dumper_1;
    df_process_monitor process_monitor_1;
    df_process_intf process_intf_2(clock,reset);
    assign process_intf_2.ap_start = AESL_inst_myproject.relu_ap_fixed_6_2_5_3_0_ap_fixed_6_2_5_3_0_relu_config3_U0.ap_start;
    assign process_intf_2.ap_ready = AESL_inst_myproject.relu_ap_fixed_6_2_5_3_0_ap_fixed_6_2_5_3_0_relu_config3_U0.ap_ready;
    assign process_intf_2.ap_done = AESL_inst_myproject.relu_ap_fixed_6_2_5_3_0_ap_fixed_6_2_5_3_0_relu_config3_U0.ap_done;
    assign process_intf_2.ap_continue = AESL_inst_myproject.relu_ap_fixed_6_2_5_3_0_ap_fixed_6_2_5_3_0_relu_config3_U0.ap_continue;
    assign process_intf_2.real_start = AESL_inst_myproject.relu_ap_fixed_6_2_5_3_0_ap_fixed_6_2_5_3_0_relu_config3_U0.ap_start;
    assign process_intf_2.pin_stall = 1'b0;
    assign process_intf_2.pout_stall = 1'b0;
    assign process_intf_2.cin_stall = 1'b0;
    assign process_intf_2.cout_stall = 1'b0;
    assign process_intf_2.region_idle = region_0_idle;
    assign process_intf_2.finish = finish;
    csv_file_dump pstall_csv_dumper_2;
    csv_file_dump pstatus_csv_dumper_2;
    df_process_monitor process_monitor_2;
    df_process_intf process_intf_3(clock,reset);
    assign process_intf_3.ap_start = AESL_inst_myproject.dense_resource_ap_fixed_6_2_5_3_0_ap_fixed_6_2_5_3_0_config5_U0.ap_start;
    assign process_intf_3.ap_ready = AESL_inst_myproject.dense_resource_ap_fixed_6_2_5_3_0_ap_fixed_6_2_5_3_0_config5_U0.ap_ready;
    assign process_intf_3.ap_done = AESL_inst_myproject.dense_resource_ap_fixed_6_2_5_3_0_ap_fixed_6_2_5_3_0_config5_U0.ap_done;
    assign process_intf_3.ap_continue = AESL_inst_myproject.dense_resource_ap_fixed_6_2_5_3_0_ap_fixed_6_2_5_3_0_config5_U0.ap_continue;
    assign process_intf_3.real_start = AESL_inst_myproject.dense_resource_ap_fixed_6_2_5_3_0_ap_fixed_6_2_5_3_0_config5_U0.ap_start;
    assign process_intf_3.pin_stall = 1'b0;
    assign process_intf_3.pout_stall = 1'b0;
    assign process_intf_3.cin_stall = 1'b0;
    assign process_intf_3.cout_stall = 1'b0;
    assign process_intf_3.region_idle = region_0_idle;
    assign process_intf_3.finish = finish;
    csv_file_dump pstall_csv_dumper_3;
    csv_file_dump pstatus_csv_dumper_3;
    df_process_monitor process_monitor_3;
    df_process_intf process_intf_4(clock,reset);
    assign process_intf_4.ap_start = AESL_inst_myproject.softmax_stable_ap_fixed_ap_fixed_6_2_5_3_0_softmax_config6_U0.ap_start;
    assign process_intf_4.ap_ready = AESL_inst_myproject.softmax_stable_ap_fixed_ap_fixed_6_2_5_3_0_softmax_config6_U0.ap_ready;
    assign process_intf_4.ap_done = AESL_inst_myproject.softmax_stable_ap_fixed_ap_fixed_6_2_5_3_0_softmax_config6_U0.ap_done;
    assign process_intf_4.ap_continue = AESL_inst_myproject.softmax_stable_ap_fixed_ap_fixed_6_2_5_3_0_softmax_config6_U0.ap_continue;
    assign process_intf_4.real_start = AESL_inst_myproject.softmax_stable_ap_fixed_ap_fixed_6_2_5_3_0_softmax_config6_U0.ap_start;
    assign process_intf_4.pin_stall = 1'b0;
    assign process_intf_4.pout_stall = 1'b0;
    assign process_intf_4.cin_stall = 1'b0;
    assign process_intf_4.cout_stall = 1'b0;
    assign process_intf_4.region_idle = region_0_idle;
    assign process_intf_4.finish = finish;
    csv_file_dump pstall_csv_dumper_4;
    csv_file_dump pstatus_csv_dumper_4;
    df_process_monitor process_monitor_4;

    nodf_module_intf module_intf_1(clock,reset);
    assign module_intf_1.ap_start = AESL_inst_myproject.ap_start;
    assign module_intf_1.ap_ready = AESL_inst_myproject.ap_ready;
    assign module_intf_1.ap_done = AESL_inst_myproject.ap_done;
    assign module_intf_1.ap_continue = 1'b1;
    assign module_intf_1.finish = finish;
    csv_file_dump mstatus_csv_dumper_1;
    nodf_module_monitor module_monitor_1;
    nodf_module_intf module_intf_2(clock,reset);
    assign module_intf_2.ap_start = 1'b0;
    assign module_intf_2.ap_ready = AESL_inst_myproject.conv_2d_cl_ap_fixed_6_2_5_3_0_ap_fixed_6_2_5_3_0_config2_U0.call_ret_fill_buffer_fu_6862.ap_ready;
    assign module_intf_2.ap_done = 1'b0;
    assign module_intf_2.ap_continue = 1'b0;
    assign module_intf_2.finish = finish;
    csv_file_dump mstatus_csv_dumper_2;
    nodf_module_monitor module_monitor_2;
    nodf_module_intf module_intf_3(clock,reset);
    assign module_intf_3.ap_start = AESL_inst_myproject.dense_resource_ap_fixed_6_2_5_3_0_ap_fixed_6_2_5_3_0_config5_U0.grp_dense_resource_rf_leq_nin_ap_fixed_ap_fixed_6_2_5_3_0_config5_s_fu_10822.ap_start;
    assign module_intf_3.ap_ready = AESL_inst_myproject.dense_resource_ap_fixed_6_2_5_3_0_ap_fixed_6_2_5_3_0_config5_U0.grp_dense_resource_rf_leq_nin_ap_fixed_ap_fixed_6_2_5_3_0_config5_s_fu_10822.ap_ready;
    assign module_intf_3.ap_done = AESL_inst_myproject.dense_resource_ap_fixed_6_2_5_3_0_ap_fixed_6_2_5_3_0_config5_U0.grp_dense_resource_rf_leq_nin_ap_fixed_ap_fixed_6_2_5_3_0_config5_s_fu_10822.ap_done;
    assign module_intf_3.ap_continue = 1'b1;
    assign module_intf_3.finish = finish;
    csv_file_dump mstatus_csv_dumper_3;
    nodf_module_monitor module_monitor_3;

    seq_loop_intf#(4) seq_loop_intf_1(clock,reset);
    assign seq_loop_intf_1.pre_loop_state0 = AESL_inst_myproject.conv_2d_cl_ap_fixed_6_2_5_3_0_ap_fixed_6_2_5_3_0_config2_U0.ap_ST_fsm_state1;
    assign seq_loop_intf_1.pre_states_valid = 1'b1;
    assign seq_loop_intf_1.post_loop_state0 = AESL_inst_myproject.conv_2d_cl_ap_fixed_6_2_5_3_0_ap_fixed_6_2_5_3_0_config2_U0.ap_ST_fsm_state4;
    assign seq_loop_intf_1.post_states_valid = 1'b1;
    assign seq_loop_intf_1.quit_loop_state0 = AESL_inst_myproject.conv_2d_cl_ap_fixed_6_2_5_3_0_ap_fixed_6_2_5_3_0_config2_U0.ap_ST_fsm_state3;
    assign seq_loop_intf_1.quit_states_valid = 1'b1;
    assign seq_loop_intf_1.cur_state = AESL_inst_myproject.conv_2d_cl_ap_fixed_6_2_5_3_0_ap_fixed_6_2_5_3_0_config2_U0.ap_CS_fsm;
    assign seq_loop_intf_1.iter_start_state = AESL_inst_myproject.conv_2d_cl_ap_fixed_6_2_5_3_0_ap_fixed_6_2_5_3_0_config2_U0.ap_ST_fsm_state2;
    assign seq_loop_intf_1.iter_end_state0 = AESL_inst_myproject.conv_2d_cl_ap_fixed_6_2_5_3_0_ap_fixed_6_2_5_3_0_config2_U0.ap_ST_fsm_state3;
    assign seq_loop_intf_1.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_1.one_state_loop = 1'b0;
    assign seq_loop_intf_1.one_state_block = 1'b0;
    assign seq_loop_intf_1.finish = finish;
    csv_file_dump seq_loop_csv_dumper_1;
    seq_loop_monitor #(4) seq_loop_monitor_1;
    upc_loop_intf#(1) upc_loop_intf_1(clock,reset);
    assign upc_loop_intf_1.cur_state = AESL_inst_myproject.dense_resource_ap_fixed_6_2_5_3_0_ap_fixed_6_2_5_3_0_config5_U0.grp_dense_resource_rf_leq_nin_ap_fixed_ap_fixed_6_2_5_3_0_config5_s_fu_10822.ap_CS_fsm;
    assign upc_loop_intf_1.iter_start_state = AESL_inst_myproject.dense_resource_ap_fixed_6_2_5_3_0_ap_fixed_6_2_5_3_0_config5_U0.grp_dense_resource_rf_leq_nin_ap_fixed_ap_fixed_6_2_5_3_0_config5_s_fu_10822.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.iter_end_state = AESL_inst_myproject.dense_resource_ap_fixed_6_2_5_3_0_ap_fixed_6_2_5_3_0_config5_U0.grp_dense_resource_rf_leq_nin_ap_fixed_ap_fixed_6_2_5_3_0_config5_s_fu_10822.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.quit_state = AESL_inst_myproject.dense_resource_ap_fixed_6_2_5_3_0_ap_fixed_6_2_5_3_0_config5_U0.grp_dense_resource_rf_leq_nin_ap_fixed_ap_fixed_6_2_5_3_0_config5_s_fu_10822.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.iter_start_block = AESL_inst_myproject.dense_resource_ap_fixed_6_2_5_3_0_ap_fixed_6_2_5_3_0_config5_U0.grp_dense_resource_rf_leq_nin_ap_fixed_ap_fixed_6_2_5_3_0_config5_s_fu_10822.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.iter_end_block = AESL_inst_myproject.dense_resource_ap_fixed_6_2_5_3_0_ap_fixed_6_2_5_3_0_config5_U0.grp_dense_resource_rf_leq_nin_ap_fixed_ap_fixed_6_2_5_3_0_config5_s_fu_10822.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.quit_block = AESL_inst_myproject.dense_resource_ap_fixed_6_2_5_3_0_ap_fixed_6_2_5_3_0_config5_U0.grp_dense_resource_rf_leq_nin_ap_fixed_ap_fixed_6_2_5_3_0_config5_s_fu_10822.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.iter_start_enable = AESL_inst_myproject.dense_resource_ap_fixed_6_2_5_3_0_ap_fixed_6_2_5_3_0_config5_U0.grp_dense_resource_rf_leq_nin_ap_fixed_ap_fixed_6_2_5_3_0_config5_s_fu_10822.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_1.iter_end_enable = AESL_inst_myproject.dense_resource_ap_fixed_6_2_5_3_0_ap_fixed_6_2_5_3_0_config5_U0.grp_dense_resource_rf_leq_nin_ap_fixed_ap_fixed_6_2_5_3_0_config5_s_fu_10822.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_1.quit_enable = AESL_inst_myproject.dense_resource_ap_fixed_6_2_5_3_0_ap_fixed_6_2_5_3_0_config5_U0.grp_dense_resource_rf_leq_nin_ap_fixed_ap_fixed_6_2_5_3_0_config5_s_fu_10822.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_1.loop_start = AESL_inst_myproject.dense_resource_ap_fixed_6_2_5_3_0_ap_fixed_6_2_5_3_0_config5_U0.grp_dense_resource_rf_leq_nin_ap_fixed_ap_fixed_6_2_5_3_0_config5_s_fu_10822.ap_start;
    assign upc_loop_intf_1.loop_ready = AESL_inst_myproject.dense_resource_ap_fixed_6_2_5_3_0_ap_fixed_6_2_5_3_0_config5_U0.grp_dense_resource_rf_leq_nin_ap_fixed_ap_fixed_6_2_5_3_0_config5_s_fu_10822.ap_ready;
    assign upc_loop_intf_1.loop_done = AESL_inst_myproject.dense_resource_ap_fixed_6_2_5_3_0_ap_fixed_6_2_5_3_0_config5_U0.grp_dense_resource_rf_leq_nin_ap_fixed_ap_fixed_6_2_5_3_0_config5_s_fu_10822.ap_done_int;
    assign upc_loop_intf_1.loop_continue = 1'b1;
    assign upc_loop_intf_1.quit_at_end = 1'b1;
    assign upc_loop_intf_1.finish = finish;
    csv_file_dump upc_loop_csv_dumper_1;
    upc_loop_monitor #(1) upc_loop_monitor_1;

    sample_manager sample_manager_inst;

initial begin
    sample_manager_inst = new;

    fifo_csv_dumper_1 = new("./depth1.csv");
    cstatus_csv_dumper_1 = new("./chan_status1.csv");
    fifo_monitor_1 = new(fifo_csv_dumper_1,fifo_intf_1,cstatus_csv_dumper_1);
    fifo_csv_dumper_2 = new("./depth2.csv");
    cstatus_csv_dumper_2 = new("./chan_status2.csv");
    fifo_monitor_2 = new(fifo_csv_dumper_2,fifo_intf_2,cstatus_csv_dumper_2);
    fifo_csv_dumper_3 = new("./depth3.csv");
    cstatus_csv_dumper_3 = new("./chan_status3.csv");
    fifo_monitor_3 = new(fifo_csv_dumper_3,fifo_intf_3,cstatus_csv_dumper_3);
    fifo_csv_dumper_4 = new("./depth4.csv");
    cstatus_csv_dumper_4 = new("./chan_status4.csv");
    fifo_monitor_4 = new(fifo_csv_dumper_4,fifo_intf_4,cstatus_csv_dumper_4);
    fifo_csv_dumper_5 = new("./depth5.csv");
    cstatus_csv_dumper_5 = new("./chan_status5.csv");
    fifo_monitor_5 = new(fifo_csv_dumper_5,fifo_intf_5,cstatus_csv_dumper_5);
    fifo_csv_dumper_6 = new("./depth6.csv");
    cstatus_csv_dumper_6 = new("./chan_status6.csv");
    fifo_monitor_6 = new(fifo_csv_dumper_6,fifo_intf_6,cstatus_csv_dumper_6);
    fifo_csv_dumper_7 = new("./depth7.csv");
    cstatus_csv_dumper_7 = new("./chan_status7.csv");
    fifo_monitor_7 = new(fifo_csv_dumper_7,fifo_intf_7,cstatus_csv_dumper_7);
    fifo_csv_dumper_8 = new("./depth8.csv");
    cstatus_csv_dumper_8 = new("./chan_status8.csv");
    fifo_monitor_8 = new(fifo_csv_dumper_8,fifo_intf_8,cstatus_csv_dumper_8);
    fifo_csv_dumper_9 = new("./depth9.csv");
    cstatus_csv_dumper_9 = new("./chan_status9.csv");
    fifo_monitor_9 = new(fifo_csv_dumper_9,fifo_intf_9,cstatus_csv_dumper_9);
    fifo_csv_dumper_10 = new("./depth10.csv");
    cstatus_csv_dumper_10 = new("./chan_status10.csv");
    fifo_monitor_10 = new(fifo_csv_dumper_10,fifo_intf_10,cstatus_csv_dumper_10);
    fifo_csv_dumper_11 = new("./depth11.csv");
    cstatus_csv_dumper_11 = new("./chan_status11.csv");
    fifo_monitor_11 = new(fifo_csv_dumper_11,fifo_intf_11,cstatus_csv_dumper_11);
    fifo_csv_dumper_12 = new("./depth12.csv");
    cstatus_csv_dumper_12 = new("./chan_status12.csv");
    fifo_monitor_12 = new(fifo_csv_dumper_12,fifo_intf_12,cstatus_csv_dumper_12);
    fifo_csv_dumper_13 = new("./depth13.csv");
    cstatus_csv_dumper_13 = new("./chan_status13.csv");
    fifo_monitor_13 = new(fifo_csv_dumper_13,fifo_intf_13,cstatus_csv_dumper_13);
    fifo_csv_dumper_14 = new("./depth14.csv");
    cstatus_csv_dumper_14 = new("./chan_status14.csv");
    fifo_monitor_14 = new(fifo_csv_dumper_14,fifo_intf_14,cstatus_csv_dumper_14);
    fifo_csv_dumper_15 = new("./depth15.csv");
    cstatus_csv_dumper_15 = new("./chan_status15.csv");
    fifo_monitor_15 = new(fifo_csv_dumper_15,fifo_intf_15,cstatus_csv_dumper_15);
    fifo_csv_dumper_16 = new("./depth16.csv");
    cstatus_csv_dumper_16 = new("./chan_status16.csv");
    fifo_monitor_16 = new(fifo_csv_dumper_16,fifo_intf_16,cstatus_csv_dumper_16);
    fifo_csv_dumper_17 = new("./depth17.csv");
    cstatus_csv_dumper_17 = new("./chan_status17.csv");
    fifo_monitor_17 = new(fifo_csv_dumper_17,fifo_intf_17,cstatus_csv_dumper_17);
    fifo_csv_dumper_18 = new("./depth18.csv");
    cstatus_csv_dumper_18 = new("./chan_status18.csv");
    fifo_monitor_18 = new(fifo_csv_dumper_18,fifo_intf_18,cstatus_csv_dumper_18);
    fifo_csv_dumper_19 = new("./depth19.csv");
    cstatus_csv_dumper_19 = new("./chan_status19.csv");
    fifo_monitor_19 = new(fifo_csv_dumper_19,fifo_intf_19,cstatus_csv_dumper_19);
    fifo_csv_dumper_20 = new("./depth20.csv");
    cstatus_csv_dumper_20 = new("./chan_status20.csv");
    fifo_monitor_20 = new(fifo_csv_dumper_20,fifo_intf_20,cstatus_csv_dumper_20);
    fifo_csv_dumper_21 = new("./depth21.csv");
    cstatus_csv_dumper_21 = new("./chan_status21.csv");
    fifo_monitor_21 = new(fifo_csv_dumper_21,fifo_intf_21,cstatus_csv_dumper_21);
    fifo_csv_dumper_22 = new("./depth22.csv");
    cstatus_csv_dumper_22 = new("./chan_status22.csv");
    fifo_monitor_22 = new(fifo_csv_dumper_22,fifo_intf_22,cstatus_csv_dumper_22);
    fifo_csv_dumper_23 = new("./depth23.csv");
    cstatus_csv_dumper_23 = new("./chan_status23.csv");
    fifo_monitor_23 = new(fifo_csv_dumper_23,fifo_intf_23,cstatus_csv_dumper_23);
    fifo_csv_dumper_24 = new("./depth24.csv");
    cstatus_csv_dumper_24 = new("./chan_status24.csv");
    fifo_monitor_24 = new(fifo_csv_dumper_24,fifo_intf_24,cstatus_csv_dumper_24);
    fifo_csv_dumper_25 = new("./depth25.csv");
    cstatus_csv_dumper_25 = new("./chan_status25.csv");
    fifo_monitor_25 = new(fifo_csv_dumper_25,fifo_intf_25,cstatus_csv_dumper_25);
    fifo_csv_dumper_26 = new("./depth26.csv");
    cstatus_csv_dumper_26 = new("./chan_status26.csv");
    fifo_monitor_26 = new(fifo_csv_dumper_26,fifo_intf_26,cstatus_csv_dumper_26);
    fifo_csv_dumper_27 = new("./depth27.csv");
    cstatus_csv_dumper_27 = new("./chan_status27.csv");
    fifo_monitor_27 = new(fifo_csv_dumper_27,fifo_intf_27,cstatus_csv_dumper_27);
    fifo_csv_dumper_28 = new("./depth28.csv");
    cstatus_csv_dumper_28 = new("./chan_status28.csv");
    fifo_monitor_28 = new(fifo_csv_dumper_28,fifo_intf_28,cstatus_csv_dumper_28);
    fifo_csv_dumper_29 = new("./depth29.csv");
    cstatus_csv_dumper_29 = new("./chan_status29.csv");
    fifo_monitor_29 = new(fifo_csv_dumper_29,fifo_intf_29,cstatus_csv_dumper_29);
    fifo_csv_dumper_30 = new("./depth30.csv");
    cstatus_csv_dumper_30 = new("./chan_status30.csv");
    fifo_monitor_30 = new(fifo_csv_dumper_30,fifo_intf_30,cstatus_csv_dumper_30);
    fifo_csv_dumper_31 = new("./depth31.csv");
    cstatus_csv_dumper_31 = new("./chan_status31.csv");
    fifo_monitor_31 = new(fifo_csv_dumper_31,fifo_intf_31,cstatus_csv_dumper_31);
    fifo_csv_dumper_32 = new("./depth32.csv");
    cstatus_csv_dumper_32 = new("./chan_status32.csv");
    fifo_monitor_32 = new(fifo_csv_dumper_32,fifo_intf_32,cstatus_csv_dumper_32);
    fifo_csv_dumper_33 = new("./depth33.csv");
    cstatus_csv_dumper_33 = new("./chan_status33.csv");
    fifo_monitor_33 = new(fifo_csv_dumper_33,fifo_intf_33,cstatus_csv_dumper_33);
    fifo_csv_dumper_34 = new("./depth34.csv");
    cstatus_csv_dumper_34 = new("./chan_status34.csv");
    fifo_monitor_34 = new(fifo_csv_dumper_34,fifo_intf_34,cstatus_csv_dumper_34);
    fifo_csv_dumper_35 = new("./depth35.csv");
    cstatus_csv_dumper_35 = new("./chan_status35.csv");
    fifo_monitor_35 = new(fifo_csv_dumper_35,fifo_intf_35,cstatus_csv_dumper_35);
    fifo_csv_dumper_36 = new("./depth36.csv");
    cstatus_csv_dumper_36 = new("./chan_status36.csv");
    fifo_monitor_36 = new(fifo_csv_dumper_36,fifo_intf_36,cstatus_csv_dumper_36);
    fifo_csv_dumper_37 = new("./depth37.csv");
    cstatus_csv_dumper_37 = new("./chan_status37.csv");
    fifo_monitor_37 = new(fifo_csv_dumper_37,fifo_intf_37,cstatus_csv_dumper_37);
    fifo_csv_dumper_38 = new("./depth38.csv");
    cstatus_csv_dumper_38 = new("./chan_status38.csv");
    fifo_monitor_38 = new(fifo_csv_dumper_38,fifo_intf_38,cstatus_csv_dumper_38);
    fifo_csv_dumper_39 = new("./depth39.csv");
    cstatus_csv_dumper_39 = new("./chan_status39.csv");
    fifo_monitor_39 = new(fifo_csv_dumper_39,fifo_intf_39,cstatus_csv_dumper_39);
    fifo_csv_dumper_40 = new("./depth40.csv");
    cstatus_csv_dumper_40 = new("./chan_status40.csv");
    fifo_monitor_40 = new(fifo_csv_dumper_40,fifo_intf_40,cstatus_csv_dumper_40);
    fifo_csv_dumper_41 = new("./depth41.csv");
    cstatus_csv_dumper_41 = new("./chan_status41.csv");
    fifo_monitor_41 = new(fifo_csv_dumper_41,fifo_intf_41,cstatus_csv_dumper_41);
    fifo_csv_dumper_42 = new("./depth42.csv");
    cstatus_csv_dumper_42 = new("./chan_status42.csv");
    fifo_monitor_42 = new(fifo_csv_dumper_42,fifo_intf_42,cstatus_csv_dumper_42);
    fifo_csv_dumper_43 = new("./depth43.csv");
    cstatus_csv_dumper_43 = new("./chan_status43.csv");
    fifo_monitor_43 = new(fifo_csv_dumper_43,fifo_intf_43,cstatus_csv_dumper_43);
    fifo_csv_dumper_44 = new("./depth44.csv");
    cstatus_csv_dumper_44 = new("./chan_status44.csv");
    fifo_monitor_44 = new(fifo_csv_dumper_44,fifo_intf_44,cstatus_csv_dumper_44);
    fifo_csv_dumper_45 = new("./depth45.csv");
    cstatus_csv_dumper_45 = new("./chan_status45.csv");
    fifo_monitor_45 = new(fifo_csv_dumper_45,fifo_intf_45,cstatus_csv_dumper_45);
    fifo_csv_dumper_46 = new("./depth46.csv");
    cstatus_csv_dumper_46 = new("./chan_status46.csv");
    fifo_monitor_46 = new(fifo_csv_dumper_46,fifo_intf_46,cstatus_csv_dumper_46);
    fifo_csv_dumper_47 = new("./depth47.csv");
    cstatus_csv_dumper_47 = new("./chan_status47.csv");
    fifo_monitor_47 = new(fifo_csv_dumper_47,fifo_intf_47,cstatus_csv_dumper_47);
    fifo_csv_dumper_48 = new("./depth48.csv");
    cstatus_csv_dumper_48 = new("./chan_status48.csv");
    fifo_monitor_48 = new(fifo_csv_dumper_48,fifo_intf_48,cstatus_csv_dumper_48);
    fifo_csv_dumper_49 = new("./depth49.csv");
    cstatus_csv_dumper_49 = new("./chan_status49.csv");
    fifo_monitor_49 = new(fifo_csv_dumper_49,fifo_intf_49,cstatus_csv_dumper_49);
    fifo_csv_dumper_50 = new("./depth50.csv");
    cstatus_csv_dumper_50 = new("./chan_status50.csv");
    fifo_monitor_50 = new(fifo_csv_dumper_50,fifo_intf_50,cstatus_csv_dumper_50);
    fifo_csv_dumper_51 = new("./depth51.csv");
    cstatus_csv_dumper_51 = new("./chan_status51.csv");
    fifo_monitor_51 = new(fifo_csv_dumper_51,fifo_intf_51,cstatus_csv_dumper_51);
    fifo_csv_dumper_52 = new("./depth52.csv");
    cstatus_csv_dumper_52 = new("./chan_status52.csv");
    fifo_monitor_52 = new(fifo_csv_dumper_52,fifo_intf_52,cstatus_csv_dumper_52);
    fifo_csv_dumper_53 = new("./depth53.csv");
    cstatus_csv_dumper_53 = new("./chan_status53.csv");
    fifo_monitor_53 = new(fifo_csv_dumper_53,fifo_intf_53,cstatus_csv_dumper_53);
    fifo_csv_dumper_54 = new("./depth54.csv");
    cstatus_csv_dumper_54 = new("./chan_status54.csv");
    fifo_monitor_54 = new(fifo_csv_dumper_54,fifo_intf_54,cstatus_csv_dumper_54);
    fifo_csv_dumper_55 = new("./depth55.csv");
    cstatus_csv_dumper_55 = new("./chan_status55.csv");
    fifo_monitor_55 = new(fifo_csv_dumper_55,fifo_intf_55,cstatus_csv_dumper_55);
    fifo_csv_dumper_56 = new("./depth56.csv");
    cstatus_csv_dumper_56 = new("./chan_status56.csv");
    fifo_monitor_56 = new(fifo_csv_dumper_56,fifo_intf_56,cstatus_csv_dumper_56);
    fifo_csv_dumper_57 = new("./depth57.csv");
    cstatus_csv_dumper_57 = new("./chan_status57.csv");
    fifo_monitor_57 = new(fifo_csv_dumper_57,fifo_intf_57,cstatus_csv_dumper_57);
    fifo_csv_dumper_58 = new("./depth58.csv");
    cstatus_csv_dumper_58 = new("./chan_status58.csv");
    fifo_monitor_58 = new(fifo_csv_dumper_58,fifo_intf_58,cstatus_csv_dumper_58);
    fifo_csv_dumper_59 = new("./depth59.csv");
    cstatus_csv_dumper_59 = new("./chan_status59.csv");
    fifo_monitor_59 = new(fifo_csv_dumper_59,fifo_intf_59,cstatus_csv_dumper_59);
    fifo_csv_dumper_60 = new("./depth60.csv");
    cstatus_csv_dumper_60 = new("./chan_status60.csv");
    fifo_monitor_60 = new(fifo_csv_dumper_60,fifo_intf_60,cstatus_csv_dumper_60);
    fifo_csv_dumper_61 = new("./depth61.csv");
    cstatus_csv_dumper_61 = new("./chan_status61.csv");
    fifo_monitor_61 = new(fifo_csv_dumper_61,fifo_intf_61,cstatus_csv_dumper_61);
    fifo_csv_dumper_62 = new("./depth62.csv");
    cstatus_csv_dumper_62 = new("./chan_status62.csv");
    fifo_monitor_62 = new(fifo_csv_dumper_62,fifo_intf_62,cstatus_csv_dumper_62);
    fifo_csv_dumper_63 = new("./depth63.csv");
    cstatus_csv_dumper_63 = new("./chan_status63.csv");
    fifo_monitor_63 = new(fifo_csv_dumper_63,fifo_intf_63,cstatus_csv_dumper_63);
    fifo_csv_dumper_64 = new("./depth64.csv");
    cstatus_csv_dumper_64 = new("./chan_status64.csv");
    fifo_monitor_64 = new(fifo_csv_dumper_64,fifo_intf_64,cstatus_csv_dumper_64);
    fifo_csv_dumper_65 = new("./depth65.csv");
    cstatus_csv_dumper_65 = new("./chan_status65.csv");
    fifo_monitor_65 = new(fifo_csv_dumper_65,fifo_intf_65,cstatus_csv_dumper_65);
    fifo_csv_dumper_66 = new("./depth66.csv");
    cstatus_csv_dumper_66 = new("./chan_status66.csv");
    fifo_monitor_66 = new(fifo_csv_dumper_66,fifo_intf_66,cstatus_csv_dumper_66);
    fifo_csv_dumper_67 = new("./depth67.csv");
    cstatus_csv_dumper_67 = new("./chan_status67.csv");
    fifo_monitor_67 = new(fifo_csv_dumper_67,fifo_intf_67,cstatus_csv_dumper_67);
    fifo_csv_dumper_68 = new("./depth68.csv");
    cstatus_csv_dumper_68 = new("./chan_status68.csv");
    fifo_monitor_68 = new(fifo_csv_dumper_68,fifo_intf_68,cstatus_csv_dumper_68);
    fifo_csv_dumper_69 = new("./depth69.csv");
    cstatus_csv_dumper_69 = new("./chan_status69.csv");
    fifo_monitor_69 = new(fifo_csv_dumper_69,fifo_intf_69,cstatus_csv_dumper_69);
    fifo_csv_dumper_70 = new("./depth70.csv");
    cstatus_csv_dumper_70 = new("./chan_status70.csv");
    fifo_monitor_70 = new(fifo_csv_dumper_70,fifo_intf_70,cstatus_csv_dumper_70);
    fifo_csv_dumper_71 = new("./depth71.csv");
    cstatus_csv_dumper_71 = new("./chan_status71.csv");
    fifo_monitor_71 = new(fifo_csv_dumper_71,fifo_intf_71,cstatus_csv_dumper_71);
    fifo_csv_dumper_72 = new("./depth72.csv");
    cstatus_csv_dumper_72 = new("./chan_status72.csv");
    fifo_monitor_72 = new(fifo_csv_dumper_72,fifo_intf_72,cstatus_csv_dumper_72);
    fifo_csv_dumper_73 = new("./depth73.csv");
    cstatus_csv_dumper_73 = new("./chan_status73.csv");
    fifo_monitor_73 = new(fifo_csv_dumper_73,fifo_intf_73,cstatus_csv_dumper_73);
    fifo_csv_dumper_74 = new("./depth74.csv");
    cstatus_csv_dumper_74 = new("./chan_status74.csv");
    fifo_monitor_74 = new(fifo_csv_dumper_74,fifo_intf_74,cstatus_csv_dumper_74);
    fifo_csv_dumper_75 = new("./depth75.csv");
    cstatus_csv_dumper_75 = new("./chan_status75.csv");
    fifo_monitor_75 = new(fifo_csv_dumper_75,fifo_intf_75,cstatus_csv_dumper_75);
    fifo_csv_dumper_76 = new("./depth76.csv");
    cstatus_csv_dumper_76 = new("./chan_status76.csv");
    fifo_monitor_76 = new(fifo_csv_dumper_76,fifo_intf_76,cstatus_csv_dumper_76);
    fifo_csv_dumper_77 = new("./depth77.csv");
    cstatus_csv_dumper_77 = new("./chan_status77.csv");
    fifo_monitor_77 = new(fifo_csv_dumper_77,fifo_intf_77,cstatus_csv_dumper_77);
    fifo_csv_dumper_78 = new("./depth78.csv");
    cstatus_csv_dumper_78 = new("./chan_status78.csv");
    fifo_monitor_78 = new(fifo_csv_dumper_78,fifo_intf_78,cstatus_csv_dumper_78);
    fifo_csv_dumper_79 = new("./depth79.csv");
    cstatus_csv_dumper_79 = new("./chan_status79.csv");
    fifo_monitor_79 = new(fifo_csv_dumper_79,fifo_intf_79,cstatus_csv_dumper_79);
    fifo_csv_dumper_80 = new("./depth80.csv");
    cstatus_csv_dumper_80 = new("./chan_status80.csv");
    fifo_monitor_80 = new(fifo_csv_dumper_80,fifo_intf_80,cstatus_csv_dumper_80);
    fifo_csv_dumper_81 = new("./depth81.csv");
    cstatus_csv_dumper_81 = new("./chan_status81.csv");
    fifo_monitor_81 = new(fifo_csv_dumper_81,fifo_intf_81,cstatus_csv_dumper_81);
    fifo_csv_dumper_82 = new("./depth82.csv");
    cstatus_csv_dumper_82 = new("./chan_status82.csv");
    fifo_monitor_82 = new(fifo_csv_dumper_82,fifo_intf_82,cstatus_csv_dumper_82);
    fifo_csv_dumper_83 = new("./depth83.csv");
    cstatus_csv_dumper_83 = new("./chan_status83.csv");
    fifo_monitor_83 = new(fifo_csv_dumper_83,fifo_intf_83,cstatus_csv_dumper_83);
    fifo_csv_dumper_84 = new("./depth84.csv");
    cstatus_csv_dumper_84 = new("./chan_status84.csv");
    fifo_monitor_84 = new(fifo_csv_dumper_84,fifo_intf_84,cstatus_csv_dumper_84);
    fifo_csv_dumper_85 = new("./depth85.csv");
    cstatus_csv_dumper_85 = new("./chan_status85.csv");
    fifo_monitor_85 = new(fifo_csv_dumper_85,fifo_intf_85,cstatus_csv_dumper_85);
    fifo_csv_dumper_86 = new("./depth86.csv");
    cstatus_csv_dumper_86 = new("./chan_status86.csv");
    fifo_monitor_86 = new(fifo_csv_dumper_86,fifo_intf_86,cstatus_csv_dumper_86);
    fifo_csv_dumper_87 = new("./depth87.csv");
    cstatus_csv_dumper_87 = new("./chan_status87.csv");
    fifo_monitor_87 = new(fifo_csv_dumper_87,fifo_intf_87,cstatus_csv_dumper_87);
    fifo_csv_dumper_88 = new("./depth88.csv");
    cstatus_csv_dumper_88 = new("./chan_status88.csv");
    fifo_monitor_88 = new(fifo_csv_dumper_88,fifo_intf_88,cstatus_csv_dumper_88);
    fifo_csv_dumper_89 = new("./depth89.csv");
    cstatus_csv_dumper_89 = new("./chan_status89.csv");
    fifo_monitor_89 = new(fifo_csv_dumper_89,fifo_intf_89,cstatus_csv_dumper_89);
    fifo_csv_dumper_90 = new("./depth90.csv");
    cstatus_csv_dumper_90 = new("./chan_status90.csv");
    fifo_monitor_90 = new(fifo_csv_dumper_90,fifo_intf_90,cstatus_csv_dumper_90);
    fifo_csv_dumper_91 = new("./depth91.csv");
    cstatus_csv_dumper_91 = new("./chan_status91.csv");
    fifo_monitor_91 = new(fifo_csv_dumper_91,fifo_intf_91,cstatus_csv_dumper_91);
    fifo_csv_dumper_92 = new("./depth92.csv");
    cstatus_csv_dumper_92 = new("./chan_status92.csv");
    fifo_monitor_92 = new(fifo_csv_dumper_92,fifo_intf_92,cstatus_csv_dumper_92);
    fifo_csv_dumper_93 = new("./depth93.csv");
    cstatus_csv_dumper_93 = new("./chan_status93.csv");
    fifo_monitor_93 = new(fifo_csv_dumper_93,fifo_intf_93,cstatus_csv_dumper_93);
    fifo_csv_dumper_94 = new("./depth94.csv");
    cstatus_csv_dumper_94 = new("./chan_status94.csv");
    fifo_monitor_94 = new(fifo_csv_dumper_94,fifo_intf_94,cstatus_csv_dumper_94);
    fifo_csv_dumper_95 = new("./depth95.csv");
    cstatus_csv_dumper_95 = new("./chan_status95.csv");
    fifo_monitor_95 = new(fifo_csv_dumper_95,fifo_intf_95,cstatus_csv_dumper_95);
    fifo_csv_dumper_96 = new("./depth96.csv");
    cstatus_csv_dumper_96 = new("./chan_status96.csv");
    fifo_monitor_96 = new(fifo_csv_dumper_96,fifo_intf_96,cstatus_csv_dumper_96);
    fifo_csv_dumper_97 = new("./depth97.csv");
    cstatus_csv_dumper_97 = new("./chan_status97.csv");
    fifo_monitor_97 = new(fifo_csv_dumper_97,fifo_intf_97,cstatus_csv_dumper_97);
    fifo_csv_dumper_98 = new("./depth98.csv");
    cstatus_csv_dumper_98 = new("./chan_status98.csv");
    fifo_monitor_98 = new(fifo_csv_dumper_98,fifo_intf_98,cstatus_csv_dumper_98);
    fifo_csv_dumper_99 = new("./depth99.csv");
    cstatus_csv_dumper_99 = new("./chan_status99.csv");
    fifo_monitor_99 = new(fifo_csv_dumper_99,fifo_intf_99,cstatus_csv_dumper_99);
    fifo_csv_dumper_100 = new("./depth100.csv");
    cstatus_csv_dumper_100 = new("./chan_status100.csv");
    fifo_monitor_100 = new(fifo_csv_dumper_100,fifo_intf_100,cstatus_csv_dumper_100);
    fifo_csv_dumper_101 = new("./depth101.csv");
    cstatus_csv_dumper_101 = new("./chan_status101.csv");
    fifo_monitor_101 = new(fifo_csv_dumper_101,fifo_intf_101,cstatus_csv_dumper_101);
    fifo_csv_dumper_102 = new("./depth102.csv");
    cstatus_csv_dumper_102 = new("./chan_status102.csv");
    fifo_monitor_102 = new(fifo_csv_dumper_102,fifo_intf_102,cstatus_csv_dumper_102);
    fifo_csv_dumper_103 = new("./depth103.csv");
    cstatus_csv_dumper_103 = new("./chan_status103.csv");
    fifo_monitor_103 = new(fifo_csv_dumper_103,fifo_intf_103,cstatus_csv_dumper_103);
    fifo_csv_dumper_104 = new("./depth104.csv");
    cstatus_csv_dumper_104 = new("./chan_status104.csv");
    fifo_monitor_104 = new(fifo_csv_dumper_104,fifo_intf_104,cstatus_csv_dumper_104);
    fifo_csv_dumper_105 = new("./depth105.csv");
    cstatus_csv_dumper_105 = new("./chan_status105.csv");
    fifo_monitor_105 = new(fifo_csv_dumper_105,fifo_intf_105,cstatus_csv_dumper_105);
    fifo_csv_dumper_106 = new("./depth106.csv");
    cstatus_csv_dumper_106 = new("./chan_status106.csv");
    fifo_monitor_106 = new(fifo_csv_dumper_106,fifo_intf_106,cstatus_csv_dumper_106);
    fifo_csv_dumper_107 = new("./depth107.csv");
    cstatus_csv_dumper_107 = new("./chan_status107.csv");
    fifo_monitor_107 = new(fifo_csv_dumper_107,fifo_intf_107,cstatus_csv_dumper_107);
    fifo_csv_dumper_108 = new("./depth108.csv");
    cstatus_csv_dumper_108 = new("./chan_status108.csv");
    fifo_monitor_108 = new(fifo_csv_dumper_108,fifo_intf_108,cstatus_csv_dumper_108);
    fifo_csv_dumper_109 = new("./depth109.csv");
    cstatus_csv_dumper_109 = new("./chan_status109.csv");
    fifo_monitor_109 = new(fifo_csv_dumper_109,fifo_intf_109,cstatus_csv_dumper_109);
    fifo_csv_dumper_110 = new("./depth110.csv");
    cstatus_csv_dumper_110 = new("./chan_status110.csv");
    fifo_monitor_110 = new(fifo_csv_dumper_110,fifo_intf_110,cstatus_csv_dumper_110);
    fifo_csv_dumper_111 = new("./depth111.csv");
    cstatus_csv_dumper_111 = new("./chan_status111.csv");
    fifo_monitor_111 = new(fifo_csv_dumper_111,fifo_intf_111,cstatus_csv_dumper_111);
    fifo_csv_dumper_112 = new("./depth112.csv");
    cstatus_csv_dumper_112 = new("./chan_status112.csv");
    fifo_monitor_112 = new(fifo_csv_dumper_112,fifo_intf_112,cstatus_csv_dumper_112);
    fifo_csv_dumper_113 = new("./depth113.csv");
    cstatus_csv_dumper_113 = new("./chan_status113.csv");
    fifo_monitor_113 = new(fifo_csv_dumper_113,fifo_intf_113,cstatus_csv_dumper_113);
    fifo_csv_dumper_114 = new("./depth114.csv");
    cstatus_csv_dumper_114 = new("./chan_status114.csv");
    fifo_monitor_114 = new(fifo_csv_dumper_114,fifo_intf_114,cstatus_csv_dumper_114);
    fifo_csv_dumper_115 = new("./depth115.csv");
    cstatus_csv_dumper_115 = new("./chan_status115.csv");
    fifo_monitor_115 = new(fifo_csv_dumper_115,fifo_intf_115,cstatus_csv_dumper_115);
    fifo_csv_dumper_116 = new("./depth116.csv");
    cstatus_csv_dumper_116 = new("./chan_status116.csv");
    fifo_monitor_116 = new(fifo_csv_dumper_116,fifo_intf_116,cstatus_csv_dumper_116);
    fifo_csv_dumper_117 = new("./depth117.csv");
    cstatus_csv_dumper_117 = new("./chan_status117.csv");
    fifo_monitor_117 = new(fifo_csv_dumper_117,fifo_intf_117,cstatus_csv_dumper_117);
    fifo_csv_dumper_118 = new("./depth118.csv");
    cstatus_csv_dumper_118 = new("./chan_status118.csv");
    fifo_monitor_118 = new(fifo_csv_dumper_118,fifo_intf_118,cstatus_csv_dumper_118);
    fifo_csv_dumper_119 = new("./depth119.csv");
    cstatus_csv_dumper_119 = new("./chan_status119.csv");
    fifo_monitor_119 = new(fifo_csv_dumper_119,fifo_intf_119,cstatus_csv_dumper_119);
    fifo_csv_dumper_120 = new("./depth120.csv");
    cstatus_csv_dumper_120 = new("./chan_status120.csv");
    fifo_monitor_120 = new(fifo_csv_dumper_120,fifo_intf_120,cstatus_csv_dumper_120);
    fifo_csv_dumper_121 = new("./depth121.csv");
    cstatus_csv_dumper_121 = new("./chan_status121.csv");
    fifo_monitor_121 = new(fifo_csv_dumper_121,fifo_intf_121,cstatus_csv_dumper_121);
    fifo_csv_dumper_122 = new("./depth122.csv");
    cstatus_csv_dumper_122 = new("./chan_status122.csv");
    fifo_monitor_122 = new(fifo_csv_dumper_122,fifo_intf_122,cstatus_csv_dumper_122);
    fifo_csv_dumper_123 = new("./depth123.csv");
    cstatus_csv_dumper_123 = new("./chan_status123.csv");
    fifo_monitor_123 = new(fifo_csv_dumper_123,fifo_intf_123,cstatus_csv_dumper_123);
    fifo_csv_dumper_124 = new("./depth124.csv");
    cstatus_csv_dumper_124 = new("./chan_status124.csv");
    fifo_monitor_124 = new(fifo_csv_dumper_124,fifo_intf_124,cstatus_csv_dumper_124);
    fifo_csv_dumper_125 = new("./depth125.csv");
    cstatus_csv_dumper_125 = new("./chan_status125.csv");
    fifo_monitor_125 = new(fifo_csv_dumper_125,fifo_intf_125,cstatus_csv_dumper_125);
    fifo_csv_dumper_126 = new("./depth126.csv");
    cstatus_csv_dumper_126 = new("./chan_status126.csv");
    fifo_monitor_126 = new(fifo_csv_dumper_126,fifo_intf_126,cstatus_csv_dumper_126);
    fifo_csv_dumper_127 = new("./depth127.csv");
    cstatus_csv_dumper_127 = new("./chan_status127.csv");
    fifo_monitor_127 = new(fifo_csv_dumper_127,fifo_intf_127,cstatus_csv_dumper_127);
    fifo_csv_dumper_128 = new("./depth128.csv");
    cstatus_csv_dumper_128 = new("./chan_status128.csv");
    fifo_monitor_128 = new(fifo_csv_dumper_128,fifo_intf_128,cstatus_csv_dumper_128);
    fifo_csv_dumper_129 = new("./depth129.csv");
    cstatus_csv_dumper_129 = new("./chan_status129.csv");
    fifo_monitor_129 = new(fifo_csv_dumper_129,fifo_intf_129,cstatus_csv_dumper_129);
    fifo_csv_dumper_130 = new("./depth130.csv");
    cstatus_csv_dumper_130 = new("./chan_status130.csv");
    fifo_monitor_130 = new(fifo_csv_dumper_130,fifo_intf_130,cstatus_csv_dumper_130);
    fifo_csv_dumper_131 = new("./depth131.csv");
    cstatus_csv_dumper_131 = new("./chan_status131.csv");
    fifo_monitor_131 = new(fifo_csv_dumper_131,fifo_intf_131,cstatus_csv_dumper_131);
    fifo_csv_dumper_132 = new("./depth132.csv");
    cstatus_csv_dumper_132 = new("./chan_status132.csv");
    fifo_monitor_132 = new(fifo_csv_dumper_132,fifo_intf_132,cstatus_csv_dumper_132);
    fifo_csv_dumper_133 = new("./depth133.csv");
    cstatus_csv_dumper_133 = new("./chan_status133.csv");
    fifo_monitor_133 = new(fifo_csv_dumper_133,fifo_intf_133,cstatus_csv_dumper_133);
    fifo_csv_dumper_134 = new("./depth134.csv");
    cstatus_csv_dumper_134 = new("./chan_status134.csv");
    fifo_monitor_134 = new(fifo_csv_dumper_134,fifo_intf_134,cstatus_csv_dumper_134);
    fifo_csv_dumper_135 = new("./depth135.csv");
    cstatus_csv_dumper_135 = new("./chan_status135.csv");
    fifo_monitor_135 = new(fifo_csv_dumper_135,fifo_intf_135,cstatus_csv_dumper_135);
    fifo_csv_dumper_136 = new("./depth136.csv");
    cstatus_csv_dumper_136 = new("./chan_status136.csv");
    fifo_monitor_136 = new(fifo_csv_dumper_136,fifo_intf_136,cstatus_csv_dumper_136);
    fifo_csv_dumper_137 = new("./depth137.csv");
    cstatus_csv_dumper_137 = new("./chan_status137.csv");
    fifo_monitor_137 = new(fifo_csv_dumper_137,fifo_intf_137,cstatus_csv_dumper_137);
    fifo_csv_dumper_138 = new("./depth138.csv");
    cstatus_csv_dumper_138 = new("./chan_status138.csv");
    fifo_monitor_138 = new(fifo_csv_dumper_138,fifo_intf_138,cstatus_csv_dumper_138);
    fifo_csv_dumper_139 = new("./depth139.csv");
    cstatus_csv_dumper_139 = new("./chan_status139.csv");
    fifo_monitor_139 = new(fifo_csv_dumper_139,fifo_intf_139,cstatus_csv_dumper_139);
    fifo_csv_dumper_140 = new("./depth140.csv");
    cstatus_csv_dumper_140 = new("./chan_status140.csv");
    fifo_monitor_140 = new(fifo_csv_dumper_140,fifo_intf_140,cstatus_csv_dumper_140);
    fifo_csv_dumper_141 = new("./depth141.csv");
    cstatus_csv_dumper_141 = new("./chan_status141.csv");
    fifo_monitor_141 = new(fifo_csv_dumper_141,fifo_intf_141,cstatus_csv_dumper_141);
    fifo_csv_dumper_142 = new("./depth142.csv");
    cstatus_csv_dumper_142 = new("./chan_status142.csv");
    fifo_monitor_142 = new(fifo_csv_dumper_142,fifo_intf_142,cstatus_csv_dumper_142);
    fifo_csv_dumper_143 = new("./depth143.csv");
    cstatus_csv_dumper_143 = new("./chan_status143.csv");
    fifo_monitor_143 = new(fifo_csv_dumper_143,fifo_intf_143,cstatus_csv_dumper_143);
    fifo_csv_dumper_144 = new("./depth144.csv");
    cstatus_csv_dumper_144 = new("./chan_status144.csv");
    fifo_monitor_144 = new(fifo_csv_dumper_144,fifo_intf_144,cstatus_csv_dumper_144);
    fifo_csv_dumper_145 = new("./depth145.csv");
    cstatus_csv_dumper_145 = new("./chan_status145.csv");
    fifo_monitor_145 = new(fifo_csv_dumper_145,fifo_intf_145,cstatus_csv_dumper_145);
    fifo_csv_dumper_146 = new("./depth146.csv");
    cstatus_csv_dumper_146 = new("./chan_status146.csv");
    fifo_monitor_146 = new(fifo_csv_dumper_146,fifo_intf_146,cstatus_csv_dumper_146);
    fifo_csv_dumper_147 = new("./depth147.csv");
    cstatus_csv_dumper_147 = new("./chan_status147.csv");
    fifo_monitor_147 = new(fifo_csv_dumper_147,fifo_intf_147,cstatus_csv_dumper_147);
    fifo_csv_dumper_148 = new("./depth148.csv");
    cstatus_csv_dumper_148 = new("./chan_status148.csv");
    fifo_monitor_148 = new(fifo_csv_dumper_148,fifo_intf_148,cstatus_csv_dumper_148);
    fifo_csv_dumper_149 = new("./depth149.csv");
    cstatus_csv_dumper_149 = new("./chan_status149.csv");
    fifo_monitor_149 = new(fifo_csv_dumper_149,fifo_intf_149,cstatus_csv_dumper_149);
    fifo_csv_dumper_150 = new("./depth150.csv");
    cstatus_csv_dumper_150 = new("./chan_status150.csv");
    fifo_monitor_150 = new(fifo_csv_dumper_150,fifo_intf_150,cstatus_csv_dumper_150);
    fifo_csv_dumper_151 = new("./depth151.csv");
    cstatus_csv_dumper_151 = new("./chan_status151.csv");
    fifo_monitor_151 = new(fifo_csv_dumper_151,fifo_intf_151,cstatus_csv_dumper_151);
    fifo_csv_dumper_152 = new("./depth152.csv");
    cstatus_csv_dumper_152 = new("./chan_status152.csv");
    fifo_monitor_152 = new(fifo_csv_dumper_152,fifo_intf_152,cstatus_csv_dumper_152);
    fifo_csv_dumper_153 = new("./depth153.csv");
    cstatus_csv_dumper_153 = new("./chan_status153.csv");
    fifo_monitor_153 = new(fifo_csv_dumper_153,fifo_intf_153,cstatus_csv_dumper_153);
    fifo_csv_dumper_154 = new("./depth154.csv");
    cstatus_csv_dumper_154 = new("./chan_status154.csv");
    fifo_monitor_154 = new(fifo_csv_dumper_154,fifo_intf_154,cstatus_csv_dumper_154);
    fifo_csv_dumper_155 = new("./depth155.csv");
    cstatus_csv_dumper_155 = new("./chan_status155.csv");
    fifo_monitor_155 = new(fifo_csv_dumper_155,fifo_intf_155,cstatus_csv_dumper_155);
    fifo_csv_dumper_156 = new("./depth156.csv");
    cstatus_csv_dumper_156 = new("./chan_status156.csv");
    fifo_monitor_156 = new(fifo_csv_dumper_156,fifo_intf_156,cstatus_csv_dumper_156);
    fifo_csv_dumper_157 = new("./depth157.csv");
    cstatus_csv_dumper_157 = new("./chan_status157.csv");
    fifo_monitor_157 = new(fifo_csv_dumper_157,fifo_intf_157,cstatus_csv_dumper_157);
    fifo_csv_dumper_158 = new("./depth158.csv");
    cstatus_csv_dumper_158 = new("./chan_status158.csv");
    fifo_monitor_158 = new(fifo_csv_dumper_158,fifo_intf_158,cstatus_csv_dumper_158);
    fifo_csv_dumper_159 = new("./depth159.csv");
    cstatus_csv_dumper_159 = new("./chan_status159.csv");
    fifo_monitor_159 = new(fifo_csv_dumper_159,fifo_intf_159,cstatus_csv_dumper_159);
    fifo_csv_dumper_160 = new("./depth160.csv");
    cstatus_csv_dumper_160 = new("./chan_status160.csv");
    fifo_monitor_160 = new(fifo_csv_dumper_160,fifo_intf_160,cstatus_csv_dumper_160);
    fifo_csv_dumper_161 = new("./depth161.csv");
    cstatus_csv_dumper_161 = new("./chan_status161.csv");
    fifo_monitor_161 = new(fifo_csv_dumper_161,fifo_intf_161,cstatus_csv_dumper_161);
    fifo_csv_dumper_162 = new("./depth162.csv");
    cstatus_csv_dumper_162 = new("./chan_status162.csv");
    fifo_monitor_162 = new(fifo_csv_dumper_162,fifo_intf_162,cstatus_csv_dumper_162);
    fifo_csv_dumper_163 = new("./depth163.csv");
    cstatus_csv_dumper_163 = new("./chan_status163.csv");
    fifo_monitor_163 = new(fifo_csv_dumper_163,fifo_intf_163,cstatus_csv_dumper_163);
    fifo_csv_dumper_164 = new("./depth164.csv");
    cstatus_csv_dumper_164 = new("./chan_status164.csv");
    fifo_monitor_164 = new(fifo_csv_dumper_164,fifo_intf_164,cstatus_csv_dumper_164);
    fifo_csv_dumper_165 = new("./depth165.csv");
    cstatus_csv_dumper_165 = new("./chan_status165.csv");
    fifo_monitor_165 = new(fifo_csv_dumper_165,fifo_intf_165,cstatus_csv_dumper_165);
    fifo_csv_dumper_166 = new("./depth166.csv");
    cstatus_csv_dumper_166 = new("./chan_status166.csv");
    fifo_monitor_166 = new(fifo_csv_dumper_166,fifo_intf_166,cstatus_csv_dumper_166);
    fifo_csv_dumper_167 = new("./depth167.csv");
    cstatus_csv_dumper_167 = new("./chan_status167.csv");
    fifo_monitor_167 = new(fifo_csv_dumper_167,fifo_intf_167,cstatus_csv_dumper_167);
    fifo_csv_dumper_168 = new("./depth168.csv");
    cstatus_csv_dumper_168 = new("./chan_status168.csv");
    fifo_monitor_168 = new(fifo_csv_dumper_168,fifo_intf_168,cstatus_csv_dumper_168);
    fifo_csv_dumper_169 = new("./depth169.csv");
    cstatus_csv_dumper_169 = new("./chan_status169.csv");
    fifo_monitor_169 = new(fifo_csv_dumper_169,fifo_intf_169,cstatus_csv_dumper_169);
    fifo_csv_dumper_170 = new("./depth170.csv");
    cstatus_csv_dumper_170 = new("./chan_status170.csv");
    fifo_monitor_170 = new(fifo_csv_dumper_170,fifo_intf_170,cstatus_csv_dumper_170);
    fifo_csv_dumper_171 = new("./depth171.csv");
    cstatus_csv_dumper_171 = new("./chan_status171.csv");
    fifo_monitor_171 = new(fifo_csv_dumper_171,fifo_intf_171,cstatus_csv_dumper_171);
    fifo_csv_dumper_172 = new("./depth172.csv");
    cstatus_csv_dumper_172 = new("./chan_status172.csv");
    fifo_monitor_172 = new(fifo_csv_dumper_172,fifo_intf_172,cstatus_csv_dumper_172);
    fifo_csv_dumper_173 = new("./depth173.csv");
    cstatus_csv_dumper_173 = new("./chan_status173.csv");
    fifo_monitor_173 = new(fifo_csv_dumper_173,fifo_intf_173,cstatus_csv_dumper_173);
    fifo_csv_dumper_174 = new("./depth174.csv");
    cstatus_csv_dumper_174 = new("./chan_status174.csv");
    fifo_monitor_174 = new(fifo_csv_dumper_174,fifo_intf_174,cstatus_csv_dumper_174);
    fifo_csv_dumper_175 = new("./depth175.csv");
    cstatus_csv_dumper_175 = new("./chan_status175.csv");
    fifo_monitor_175 = new(fifo_csv_dumper_175,fifo_intf_175,cstatus_csv_dumper_175);
    fifo_csv_dumper_176 = new("./depth176.csv");
    cstatus_csv_dumper_176 = new("./chan_status176.csv");
    fifo_monitor_176 = new(fifo_csv_dumper_176,fifo_intf_176,cstatus_csv_dumper_176);
    fifo_csv_dumper_177 = new("./depth177.csv");
    cstatus_csv_dumper_177 = new("./chan_status177.csv");
    fifo_monitor_177 = new(fifo_csv_dumper_177,fifo_intf_177,cstatus_csv_dumper_177);
    fifo_csv_dumper_178 = new("./depth178.csv");
    cstatus_csv_dumper_178 = new("./chan_status178.csv");
    fifo_monitor_178 = new(fifo_csv_dumper_178,fifo_intf_178,cstatus_csv_dumper_178);
    fifo_csv_dumper_179 = new("./depth179.csv");
    cstatus_csv_dumper_179 = new("./chan_status179.csv");
    fifo_monitor_179 = new(fifo_csv_dumper_179,fifo_intf_179,cstatus_csv_dumper_179);
    fifo_csv_dumper_180 = new("./depth180.csv");
    cstatus_csv_dumper_180 = new("./chan_status180.csv");
    fifo_monitor_180 = new(fifo_csv_dumper_180,fifo_intf_180,cstatus_csv_dumper_180);
    fifo_csv_dumper_181 = new("./depth181.csv");
    cstatus_csv_dumper_181 = new("./chan_status181.csv");
    fifo_monitor_181 = new(fifo_csv_dumper_181,fifo_intf_181,cstatus_csv_dumper_181);
    fifo_csv_dumper_182 = new("./depth182.csv");
    cstatus_csv_dumper_182 = new("./chan_status182.csv");
    fifo_monitor_182 = new(fifo_csv_dumper_182,fifo_intf_182,cstatus_csv_dumper_182);
    fifo_csv_dumper_183 = new("./depth183.csv");
    cstatus_csv_dumper_183 = new("./chan_status183.csv");
    fifo_monitor_183 = new(fifo_csv_dumper_183,fifo_intf_183,cstatus_csv_dumper_183);
    fifo_csv_dumper_184 = new("./depth184.csv");
    cstatus_csv_dumper_184 = new("./chan_status184.csv");
    fifo_monitor_184 = new(fifo_csv_dumper_184,fifo_intf_184,cstatus_csv_dumper_184);
    fifo_csv_dumper_185 = new("./depth185.csv");
    cstatus_csv_dumper_185 = new("./chan_status185.csv");
    fifo_monitor_185 = new(fifo_csv_dumper_185,fifo_intf_185,cstatus_csv_dumper_185);
    fifo_csv_dumper_186 = new("./depth186.csv");
    cstatus_csv_dumper_186 = new("./chan_status186.csv");
    fifo_monitor_186 = new(fifo_csv_dumper_186,fifo_intf_186,cstatus_csv_dumper_186);
    fifo_csv_dumper_187 = new("./depth187.csv");
    cstatus_csv_dumper_187 = new("./chan_status187.csv");
    fifo_monitor_187 = new(fifo_csv_dumper_187,fifo_intf_187,cstatus_csv_dumper_187);
    fifo_csv_dumper_188 = new("./depth188.csv");
    cstatus_csv_dumper_188 = new("./chan_status188.csv");
    fifo_monitor_188 = new(fifo_csv_dumper_188,fifo_intf_188,cstatus_csv_dumper_188);
    fifo_csv_dumper_189 = new("./depth189.csv");
    cstatus_csv_dumper_189 = new("./chan_status189.csv");
    fifo_monitor_189 = new(fifo_csv_dumper_189,fifo_intf_189,cstatus_csv_dumper_189);
    fifo_csv_dumper_190 = new("./depth190.csv");
    cstatus_csv_dumper_190 = new("./chan_status190.csv");
    fifo_monitor_190 = new(fifo_csv_dumper_190,fifo_intf_190,cstatus_csv_dumper_190);
    fifo_csv_dumper_191 = new("./depth191.csv");
    cstatus_csv_dumper_191 = new("./chan_status191.csv");
    fifo_monitor_191 = new(fifo_csv_dumper_191,fifo_intf_191,cstatus_csv_dumper_191);
    fifo_csv_dumper_192 = new("./depth192.csv");
    cstatus_csv_dumper_192 = new("./chan_status192.csv");
    fifo_monitor_192 = new(fifo_csv_dumper_192,fifo_intf_192,cstatus_csv_dumper_192);
    fifo_csv_dumper_193 = new("./depth193.csv");
    cstatus_csv_dumper_193 = new("./chan_status193.csv");
    fifo_monitor_193 = new(fifo_csv_dumper_193,fifo_intf_193,cstatus_csv_dumper_193);
    fifo_csv_dumper_194 = new("./depth194.csv");
    cstatus_csv_dumper_194 = new("./chan_status194.csv");
    fifo_monitor_194 = new(fifo_csv_dumper_194,fifo_intf_194,cstatus_csv_dumper_194);
    fifo_csv_dumper_195 = new("./depth195.csv");
    cstatus_csv_dumper_195 = new("./chan_status195.csv");
    fifo_monitor_195 = new(fifo_csv_dumper_195,fifo_intf_195,cstatus_csv_dumper_195);
    fifo_csv_dumper_196 = new("./depth196.csv");
    cstatus_csv_dumper_196 = new("./chan_status196.csv");
    fifo_monitor_196 = new(fifo_csv_dumper_196,fifo_intf_196,cstatus_csv_dumper_196);
    fifo_csv_dumper_197 = new("./depth197.csv");
    cstatus_csv_dumper_197 = new("./chan_status197.csv");
    fifo_monitor_197 = new(fifo_csv_dumper_197,fifo_intf_197,cstatus_csv_dumper_197);
    fifo_csv_dumper_198 = new("./depth198.csv");
    cstatus_csv_dumper_198 = new("./chan_status198.csv");
    fifo_monitor_198 = new(fifo_csv_dumper_198,fifo_intf_198,cstatus_csv_dumper_198);
    fifo_csv_dumper_199 = new("./depth199.csv");
    cstatus_csv_dumper_199 = new("./chan_status199.csv");
    fifo_monitor_199 = new(fifo_csv_dumper_199,fifo_intf_199,cstatus_csv_dumper_199);
    fifo_csv_dumper_200 = new("./depth200.csv");
    cstatus_csv_dumper_200 = new("./chan_status200.csv");
    fifo_monitor_200 = new(fifo_csv_dumper_200,fifo_intf_200,cstatus_csv_dumper_200);
    fifo_csv_dumper_201 = new("./depth201.csv");
    cstatus_csv_dumper_201 = new("./chan_status201.csv");
    fifo_monitor_201 = new(fifo_csv_dumper_201,fifo_intf_201,cstatus_csv_dumper_201);
    fifo_csv_dumper_202 = new("./depth202.csv");
    cstatus_csv_dumper_202 = new("./chan_status202.csv");
    fifo_monitor_202 = new(fifo_csv_dumper_202,fifo_intf_202,cstatus_csv_dumper_202);
    fifo_csv_dumper_203 = new("./depth203.csv");
    cstatus_csv_dumper_203 = new("./chan_status203.csv");
    fifo_monitor_203 = new(fifo_csv_dumper_203,fifo_intf_203,cstatus_csv_dumper_203);
    fifo_csv_dumper_204 = new("./depth204.csv");
    cstatus_csv_dumper_204 = new("./chan_status204.csv");
    fifo_monitor_204 = new(fifo_csv_dumper_204,fifo_intf_204,cstatus_csv_dumper_204);
    fifo_csv_dumper_205 = new("./depth205.csv");
    cstatus_csv_dumper_205 = new("./chan_status205.csv");
    fifo_monitor_205 = new(fifo_csv_dumper_205,fifo_intf_205,cstatus_csv_dumper_205);
    fifo_csv_dumper_206 = new("./depth206.csv");
    cstatus_csv_dumper_206 = new("./chan_status206.csv");
    fifo_monitor_206 = new(fifo_csv_dumper_206,fifo_intf_206,cstatus_csv_dumper_206);
    fifo_csv_dumper_207 = new("./depth207.csv");
    cstatus_csv_dumper_207 = new("./chan_status207.csv");
    fifo_monitor_207 = new(fifo_csv_dumper_207,fifo_intf_207,cstatus_csv_dumper_207);
    fifo_csv_dumper_208 = new("./depth208.csv");
    cstatus_csv_dumper_208 = new("./chan_status208.csv");
    fifo_monitor_208 = new(fifo_csv_dumper_208,fifo_intf_208,cstatus_csv_dumper_208);
    fifo_csv_dumper_209 = new("./depth209.csv");
    cstatus_csv_dumper_209 = new("./chan_status209.csv");
    fifo_monitor_209 = new(fifo_csv_dumper_209,fifo_intf_209,cstatus_csv_dumper_209);
    fifo_csv_dumper_210 = new("./depth210.csv");
    cstatus_csv_dumper_210 = new("./chan_status210.csv");
    fifo_monitor_210 = new(fifo_csv_dumper_210,fifo_intf_210,cstatus_csv_dumper_210);
    fifo_csv_dumper_211 = new("./depth211.csv");
    cstatus_csv_dumper_211 = new("./chan_status211.csv");
    fifo_monitor_211 = new(fifo_csv_dumper_211,fifo_intf_211,cstatus_csv_dumper_211);
    fifo_csv_dumper_212 = new("./depth212.csv");
    cstatus_csv_dumper_212 = new("./chan_status212.csv");
    fifo_monitor_212 = new(fifo_csv_dumper_212,fifo_intf_212,cstatus_csv_dumper_212);
    fifo_csv_dumper_213 = new("./depth213.csv");
    cstatus_csv_dumper_213 = new("./chan_status213.csv");
    fifo_monitor_213 = new(fifo_csv_dumper_213,fifo_intf_213,cstatus_csv_dumper_213);
    fifo_csv_dumper_214 = new("./depth214.csv");
    cstatus_csv_dumper_214 = new("./chan_status214.csv");
    fifo_monitor_214 = new(fifo_csv_dumper_214,fifo_intf_214,cstatus_csv_dumper_214);
    fifo_csv_dumper_215 = new("./depth215.csv");
    cstatus_csv_dumper_215 = new("./chan_status215.csv");
    fifo_monitor_215 = new(fifo_csv_dumper_215,fifo_intf_215,cstatus_csv_dumper_215);
    fifo_csv_dumper_216 = new("./depth216.csv");
    cstatus_csv_dumper_216 = new("./chan_status216.csv");
    fifo_monitor_216 = new(fifo_csv_dumper_216,fifo_intf_216,cstatus_csv_dumper_216);
    fifo_csv_dumper_217 = new("./depth217.csv");
    cstatus_csv_dumper_217 = new("./chan_status217.csv");
    fifo_monitor_217 = new(fifo_csv_dumper_217,fifo_intf_217,cstatus_csv_dumper_217);
    fifo_csv_dumper_218 = new("./depth218.csv");
    cstatus_csv_dumper_218 = new("./chan_status218.csv");
    fifo_monitor_218 = new(fifo_csv_dumper_218,fifo_intf_218,cstatus_csv_dumper_218);
    fifo_csv_dumper_219 = new("./depth219.csv");
    cstatus_csv_dumper_219 = new("./chan_status219.csv");
    fifo_monitor_219 = new(fifo_csv_dumper_219,fifo_intf_219,cstatus_csv_dumper_219);
    fifo_csv_dumper_220 = new("./depth220.csv");
    cstatus_csv_dumper_220 = new("./chan_status220.csv");
    fifo_monitor_220 = new(fifo_csv_dumper_220,fifo_intf_220,cstatus_csv_dumper_220);
    fifo_csv_dumper_221 = new("./depth221.csv");
    cstatus_csv_dumper_221 = new("./chan_status221.csv");
    fifo_monitor_221 = new(fifo_csv_dumper_221,fifo_intf_221,cstatus_csv_dumper_221);
    fifo_csv_dumper_222 = new("./depth222.csv");
    cstatus_csv_dumper_222 = new("./chan_status222.csv");
    fifo_monitor_222 = new(fifo_csv_dumper_222,fifo_intf_222,cstatus_csv_dumper_222);
    fifo_csv_dumper_223 = new("./depth223.csv");
    cstatus_csv_dumper_223 = new("./chan_status223.csv");
    fifo_monitor_223 = new(fifo_csv_dumper_223,fifo_intf_223,cstatus_csv_dumper_223);
    fifo_csv_dumper_224 = new("./depth224.csv");
    cstatus_csv_dumper_224 = new("./chan_status224.csv");
    fifo_monitor_224 = new(fifo_csv_dumper_224,fifo_intf_224,cstatus_csv_dumper_224);
    fifo_csv_dumper_225 = new("./depth225.csv");
    cstatus_csv_dumper_225 = new("./chan_status225.csv");
    fifo_monitor_225 = new(fifo_csv_dumper_225,fifo_intf_225,cstatus_csv_dumper_225);
    fifo_csv_dumper_226 = new("./depth226.csv");
    cstatus_csv_dumper_226 = new("./chan_status226.csv");
    fifo_monitor_226 = new(fifo_csv_dumper_226,fifo_intf_226,cstatus_csv_dumper_226);
    fifo_csv_dumper_227 = new("./depth227.csv");
    cstatus_csv_dumper_227 = new("./chan_status227.csv");
    fifo_monitor_227 = new(fifo_csv_dumper_227,fifo_intf_227,cstatus_csv_dumper_227);
    fifo_csv_dumper_228 = new("./depth228.csv");
    cstatus_csv_dumper_228 = new("./chan_status228.csv");
    fifo_monitor_228 = new(fifo_csv_dumper_228,fifo_intf_228,cstatus_csv_dumper_228);
    fifo_csv_dumper_229 = new("./depth229.csv");
    cstatus_csv_dumper_229 = new("./chan_status229.csv");
    fifo_monitor_229 = new(fifo_csv_dumper_229,fifo_intf_229,cstatus_csv_dumper_229);
    fifo_csv_dumper_230 = new("./depth230.csv");
    cstatus_csv_dumper_230 = new("./chan_status230.csv");
    fifo_monitor_230 = new(fifo_csv_dumper_230,fifo_intf_230,cstatus_csv_dumper_230);
    fifo_csv_dumper_231 = new("./depth231.csv");
    cstatus_csv_dumper_231 = new("./chan_status231.csv");
    fifo_monitor_231 = new(fifo_csv_dumper_231,fifo_intf_231,cstatus_csv_dumper_231);
    fifo_csv_dumper_232 = new("./depth232.csv");
    cstatus_csv_dumper_232 = new("./chan_status232.csv");
    fifo_monitor_232 = new(fifo_csv_dumper_232,fifo_intf_232,cstatus_csv_dumper_232);
    fifo_csv_dumper_233 = new("./depth233.csv");
    cstatus_csv_dumper_233 = new("./chan_status233.csv");
    fifo_monitor_233 = new(fifo_csv_dumper_233,fifo_intf_233,cstatus_csv_dumper_233);
    fifo_csv_dumper_234 = new("./depth234.csv");
    cstatus_csv_dumper_234 = new("./chan_status234.csv");
    fifo_monitor_234 = new(fifo_csv_dumper_234,fifo_intf_234,cstatus_csv_dumper_234);
    fifo_csv_dumper_235 = new("./depth235.csv");
    cstatus_csv_dumper_235 = new("./chan_status235.csv");
    fifo_monitor_235 = new(fifo_csv_dumper_235,fifo_intf_235,cstatus_csv_dumper_235);
    fifo_csv_dumper_236 = new("./depth236.csv");
    cstatus_csv_dumper_236 = new("./chan_status236.csv");
    fifo_monitor_236 = new(fifo_csv_dumper_236,fifo_intf_236,cstatus_csv_dumper_236);
    fifo_csv_dumper_237 = new("./depth237.csv");
    cstatus_csv_dumper_237 = new("./chan_status237.csv");
    fifo_monitor_237 = new(fifo_csv_dumper_237,fifo_intf_237,cstatus_csv_dumper_237);
    fifo_csv_dumper_238 = new("./depth238.csv");
    cstatus_csv_dumper_238 = new("./chan_status238.csv");
    fifo_monitor_238 = new(fifo_csv_dumper_238,fifo_intf_238,cstatus_csv_dumper_238);
    fifo_csv_dumper_239 = new("./depth239.csv");
    cstatus_csv_dumper_239 = new("./chan_status239.csv");
    fifo_monitor_239 = new(fifo_csv_dumper_239,fifo_intf_239,cstatus_csv_dumper_239);
    fifo_csv_dumper_240 = new("./depth240.csv");
    cstatus_csv_dumper_240 = new("./chan_status240.csv");
    fifo_monitor_240 = new(fifo_csv_dumper_240,fifo_intf_240,cstatus_csv_dumper_240);
    fifo_csv_dumper_241 = new("./depth241.csv");
    cstatus_csv_dumper_241 = new("./chan_status241.csv");
    fifo_monitor_241 = new(fifo_csv_dumper_241,fifo_intf_241,cstatus_csv_dumper_241);
    fifo_csv_dumper_242 = new("./depth242.csv");
    cstatus_csv_dumper_242 = new("./chan_status242.csv");
    fifo_monitor_242 = new(fifo_csv_dumper_242,fifo_intf_242,cstatus_csv_dumper_242);
    fifo_csv_dumper_243 = new("./depth243.csv");
    cstatus_csv_dumper_243 = new("./chan_status243.csv");
    fifo_monitor_243 = new(fifo_csv_dumper_243,fifo_intf_243,cstatus_csv_dumper_243);
    fifo_csv_dumper_244 = new("./depth244.csv");
    cstatus_csv_dumper_244 = new("./chan_status244.csv");
    fifo_monitor_244 = new(fifo_csv_dumper_244,fifo_intf_244,cstatus_csv_dumper_244);
    fifo_csv_dumper_245 = new("./depth245.csv");
    cstatus_csv_dumper_245 = new("./chan_status245.csv");
    fifo_monitor_245 = new(fifo_csv_dumper_245,fifo_intf_245,cstatus_csv_dumper_245);
    fifo_csv_dumper_246 = new("./depth246.csv");
    cstatus_csv_dumper_246 = new("./chan_status246.csv");
    fifo_monitor_246 = new(fifo_csv_dumper_246,fifo_intf_246,cstatus_csv_dumper_246);
    fifo_csv_dumper_247 = new("./depth247.csv");
    cstatus_csv_dumper_247 = new("./chan_status247.csv");
    fifo_monitor_247 = new(fifo_csv_dumper_247,fifo_intf_247,cstatus_csv_dumper_247);
    fifo_csv_dumper_248 = new("./depth248.csv");
    cstatus_csv_dumper_248 = new("./chan_status248.csv");
    fifo_monitor_248 = new(fifo_csv_dumper_248,fifo_intf_248,cstatus_csv_dumper_248);
    fifo_csv_dumper_249 = new("./depth249.csv");
    cstatus_csv_dumper_249 = new("./chan_status249.csv");
    fifo_monitor_249 = new(fifo_csv_dumper_249,fifo_intf_249,cstatus_csv_dumper_249);
    fifo_csv_dumper_250 = new("./depth250.csv");
    cstatus_csv_dumper_250 = new("./chan_status250.csv");
    fifo_monitor_250 = new(fifo_csv_dumper_250,fifo_intf_250,cstatus_csv_dumper_250);
    fifo_csv_dumper_251 = new("./depth251.csv");
    cstatus_csv_dumper_251 = new("./chan_status251.csv");
    fifo_monitor_251 = new(fifo_csv_dumper_251,fifo_intf_251,cstatus_csv_dumper_251);
    fifo_csv_dumper_252 = new("./depth252.csv");
    cstatus_csv_dumper_252 = new("./chan_status252.csv");
    fifo_monitor_252 = new(fifo_csv_dumper_252,fifo_intf_252,cstatus_csv_dumper_252);
    fifo_csv_dumper_253 = new("./depth253.csv");
    cstatus_csv_dumper_253 = new("./chan_status253.csv");
    fifo_monitor_253 = new(fifo_csv_dumper_253,fifo_intf_253,cstatus_csv_dumper_253);
    fifo_csv_dumper_254 = new("./depth254.csv");
    cstatus_csv_dumper_254 = new("./chan_status254.csv");
    fifo_monitor_254 = new(fifo_csv_dumper_254,fifo_intf_254,cstatus_csv_dumper_254);
    fifo_csv_dumper_255 = new("./depth255.csv");
    cstatus_csv_dumper_255 = new("./chan_status255.csv");
    fifo_monitor_255 = new(fifo_csv_dumper_255,fifo_intf_255,cstatus_csv_dumper_255);
    fifo_csv_dumper_256 = new("./depth256.csv");
    cstatus_csv_dumper_256 = new("./chan_status256.csv");
    fifo_monitor_256 = new(fifo_csv_dumper_256,fifo_intf_256,cstatus_csv_dumper_256);
    fifo_csv_dumper_257 = new("./depth257.csv");
    cstatus_csv_dumper_257 = new("./chan_status257.csv");
    fifo_monitor_257 = new(fifo_csv_dumper_257,fifo_intf_257,cstatus_csv_dumper_257);
    fifo_csv_dumper_258 = new("./depth258.csv");
    cstatus_csv_dumper_258 = new("./chan_status258.csv");
    fifo_monitor_258 = new(fifo_csv_dumper_258,fifo_intf_258,cstatus_csv_dumper_258);
    fifo_csv_dumper_259 = new("./depth259.csv");
    cstatus_csv_dumper_259 = new("./chan_status259.csv");
    fifo_monitor_259 = new(fifo_csv_dumper_259,fifo_intf_259,cstatus_csv_dumper_259);
    fifo_csv_dumper_260 = new("./depth260.csv");
    cstatus_csv_dumper_260 = new("./chan_status260.csv");
    fifo_monitor_260 = new(fifo_csv_dumper_260,fifo_intf_260,cstatus_csv_dumper_260);
    fifo_csv_dumper_261 = new("./depth261.csv");
    cstatus_csv_dumper_261 = new("./chan_status261.csv");
    fifo_monitor_261 = new(fifo_csv_dumper_261,fifo_intf_261,cstatus_csv_dumper_261);
    fifo_csv_dumper_262 = new("./depth262.csv");
    cstatus_csv_dumper_262 = new("./chan_status262.csv");
    fifo_monitor_262 = new(fifo_csv_dumper_262,fifo_intf_262,cstatus_csv_dumper_262);
    fifo_csv_dumper_263 = new("./depth263.csv");
    cstatus_csv_dumper_263 = new("./chan_status263.csv");
    fifo_monitor_263 = new(fifo_csv_dumper_263,fifo_intf_263,cstatus_csv_dumper_263);
    fifo_csv_dumper_264 = new("./depth264.csv");
    cstatus_csv_dumper_264 = new("./chan_status264.csv");
    fifo_monitor_264 = new(fifo_csv_dumper_264,fifo_intf_264,cstatus_csv_dumper_264);
    fifo_csv_dumper_265 = new("./depth265.csv");
    cstatus_csv_dumper_265 = new("./chan_status265.csv");
    fifo_monitor_265 = new(fifo_csv_dumper_265,fifo_intf_265,cstatus_csv_dumper_265);
    fifo_csv_dumper_266 = new("./depth266.csv");
    cstatus_csv_dumper_266 = new("./chan_status266.csv");
    fifo_monitor_266 = new(fifo_csv_dumper_266,fifo_intf_266,cstatus_csv_dumper_266);
    fifo_csv_dumper_267 = new("./depth267.csv");
    cstatus_csv_dumper_267 = new("./chan_status267.csv");
    fifo_monitor_267 = new(fifo_csv_dumper_267,fifo_intf_267,cstatus_csv_dumper_267);
    fifo_csv_dumper_268 = new("./depth268.csv");
    cstatus_csv_dumper_268 = new("./chan_status268.csv");
    fifo_monitor_268 = new(fifo_csv_dumper_268,fifo_intf_268,cstatus_csv_dumper_268);
    fifo_csv_dumper_269 = new("./depth269.csv");
    cstatus_csv_dumper_269 = new("./chan_status269.csv");
    fifo_monitor_269 = new(fifo_csv_dumper_269,fifo_intf_269,cstatus_csv_dumper_269);
    fifo_csv_dumper_270 = new("./depth270.csv");
    cstatus_csv_dumper_270 = new("./chan_status270.csv");
    fifo_monitor_270 = new(fifo_csv_dumper_270,fifo_intf_270,cstatus_csv_dumper_270);
    fifo_csv_dumper_271 = new("./depth271.csv");
    cstatus_csv_dumper_271 = new("./chan_status271.csv");
    fifo_monitor_271 = new(fifo_csv_dumper_271,fifo_intf_271,cstatus_csv_dumper_271);
    fifo_csv_dumper_272 = new("./depth272.csv");
    cstatus_csv_dumper_272 = new("./chan_status272.csv");
    fifo_monitor_272 = new(fifo_csv_dumper_272,fifo_intf_272,cstatus_csv_dumper_272);
    fifo_csv_dumper_273 = new("./depth273.csv");
    cstatus_csv_dumper_273 = new("./chan_status273.csv");
    fifo_monitor_273 = new(fifo_csv_dumper_273,fifo_intf_273,cstatus_csv_dumper_273);
    fifo_csv_dumper_274 = new("./depth274.csv");
    cstatus_csv_dumper_274 = new("./chan_status274.csv");
    fifo_monitor_274 = new(fifo_csv_dumper_274,fifo_intf_274,cstatus_csv_dumper_274);
    fifo_csv_dumper_275 = new("./depth275.csv");
    cstatus_csv_dumper_275 = new("./chan_status275.csv");
    fifo_monitor_275 = new(fifo_csv_dumper_275,fifo_intf_275,cstatus_csv_dumper_275);
    fifo_csv_dumper_276 = new("./depth276.csv");
    cstatus_csv_dumper_276 = new("./chan_status276.csv");
    fifo_monitor_276 = new(fifo_csv_dumper_276,fifo_intf_276,cstatus_csv_dumper_276);
    fifo_csv_dumper_277 = new("./depth277.csv");
    cstatus_csv_dumper_277 = new("./chan_status277.csv");
    fifo_monitor_277 = new(fifo_csv_dumper_277,fifo_intf_277,cstatus_csv_dumper_277);
    fifo_csv_dumper_278 = new("./depth278.csv");
    cstatus_csv_dumper_278 = new("./chan_status278.csv");
    fifo_monitor_278 = new(fifo_csv_dumper_278,fifo_intf_278,cstatus_csv_dumper_278);
    fifo_csv_dumper_279 = new("./depth279.csv");
    cstatus_csv_dumper_279 = new("./chan_status279.csv");
    fifo_monitor_279 = new(fifo_csv_dumper_279,fifo_intf_279,cstatus_csv_dumper_279);
    fifo_csv_dumper_280 = new("./depth280.csv");
    cstatus_csv_dumper_280 = new("./chan_status280.csv");
    fifo_monitor_280 = new(fifo_csv_dumper_280,fifo_intf_280,cstatus_csv_dumper_280);
    fifo_csv_dumper_281 = new("./depth281.csv");
    cstatus_csv_dumper_281 = new("./chan_status281.csv");
    fifo_monitor_281 = new(fifo_csv_dumper_281,fifo_intf_281,cstatus_csv_dumper_281);
    fifo_csv_dumper_282 = new("./depth282.csv");
    cstatus_csv_dumper_282 = new("./chan_status282.csv");
    fifo_monitor_282 = new(fifo_csv_dumper_282,fifo_intf_282,cstatus_csv_dumper_282);
    fifo_csv_dumper_283 = new("./depth283.csv");
    cstatus_csv_dumper_283 = new("./chan_status283.csv");
    fifo_monitor_283 = new(fifo_csv_dumper_283,fifo_intf_283,cstatus_csv_dumper_283);
    fifo_csv_dumper_284 = new("./depth284.csv");
    cstatus_csv_dumper_284 = new("./chan_status284.csv");
    fifo_monitor_284 = new(fifo_csv_dumper_284,fifo_intf_284,cstatus_csv_dumper_284);
    fifo_csv_dumper_285 = new("./depth285.csv");
    cstatus_csv_dumper_285 = new("./chan_status285.csv");
    fifo_monitor_285 = new(fifo_csv_dumper_285,fifo_intf_285,cstatus_csv_dumper_285);
    fifo_csv_dumper_286 = new("./depth286.csv");
    cstatus_csv_dumper_286 = new("./chan_status286.csv");
    fifo_monitor_286 = new(fifo_csv_dumper_286,fifo_intf_286,cstatus_csv_dumper_286);
    fifo_csv_dumper_287 = new("./depth287.csv");
    cstatus_csv_dumper_287 = new("./chan_status287.csv");
    fifo_monitor_287 = new(fifo_csv_dumper_287,fifo_intf_287,cstatus_csv_dumper_287);
    fifo_csv_dumper_288 = new("./depth288.csv");
    cstatus_csv_dumper_288 = new("./chan_status288.csv");
    fifo_monitor_288 = new(fifo_csv_dumper_288,fifo_intf_288,cstatus_csv_dumper_288);
    fifo_csv_dumper_289 = new("./depth289.csv");
    cstatus_csv_dumper_289 = new("./chan_status289.csv");
    fifo_monitor_289 = new(fifo_csv_dumper_289,fifo_intf_289,cstatus_csv_dumper_289);
    fifo_csv_dumper_290 = new("./depth290.csv");
    cstatus_csv_dumper_290 = new("./chan_status290.csv");
    fifo_monitor_290 = new(fifo_csv_dumper_290,fifo_intf_290,cstatus_csv_dumper_290);
    fifo_csv_dumper_291 = new("./depth291.csv");
    cstatus_csv_dumper_291 = new("./chan_status291.csv");
    fifo_monitor_291 = new(fifo_csv_dumper_291,fifo_intf_291,cstatus_csv_dumper_291);
    fifo_csv_dumper_292 = new("./depth292.csv");
    cstatus_csv_dumper_292 = new("./chan_status292.csv");
    fifo_monitor_292 = new(fifo_csv_dumper_292,fifo_intf_292,cstatus_csv_dumper_292);
    fifo_csv_dumper_293 = new("./depth293.csv");
    cstatus_csv_dumper_293 = new("./chan_status293.csv");
    fifo_monitor_293 = new(fifo_csv_dumper_293,fifo_intf_293,cstatus_csv_dumper_293);
    fifo_csv_dumper_294 = new("./depth294.csv");
    cstatus_csv_dumper_294 = new("./chan_status294.csv");
    fifo_monitor_294 = new(fifo_csv_dumper_294,fifo_intf_294,cstatus_csv_dumper_294);
    fifo_csv_dumper_295 = new("./depth295.csv");
    cstatus_csv_dumper_295 = new("./chan_status295.csv");
    fifo_monitor_295 = new(fifo_csv_dumper_295,fifo_intf_295,cstatus_csv_dumper_295);
    fifo_csv_dumper_296 = new("./depth296.csv");
    cstatus_csv_dumper_296 = new("./chan_status296.csv");
    fifo_monitor_296 = new(fifo_csv_dumper_296,fifo_intf_296,cstatus_csv_dumper_296);
    fifo_csv_dumper_297 = new("./depth297.csv");
    cstatus_csv_dumper_297 = new("./chan_status297.csv");
    fifo_monitor_297 = new(fifo_csv_dumper_297,fifo_intf_297,cstatus_csv_dumper_297);
    fifo_csv_dumper_298 = new("./depth298.csv");
    cstatus_csv_dumper_298 = new("./chan_status298.csv");
    fifo_monitor_298 = new(fifo_csv_dumper_298,fifo_intf_298,cstatus_csv_dumper_298);
    fifo_csv_dumper_299 = new("./depth299.csv");
    cstatus_csv_dumper_299 = new("./chan_status299.csv");
    fifo_monitor_299 = new(fifo_csv_dumper_299,fifo_intf_299,cstatus_csv_dumper_299);
    fifo_csv_dumper_300 = new("./depth300.csv");
    cstatus_csv_dumper_300 = new("./chan_status300.csv");
    fifo_monitor_300 = new(fifo_csv_dumper_300,fifo_intf_300,cstatus_csv_dumper_300);
    fifo_csv_dumper_301 = new("./depth301.csv");
    cstatus_csv_dumper_301 = new("./chan_status301.csv");
    fifo_monitor_301 = new(fifo_csv_dumper_301,fifo_intf_301,cstatus_csv_dumper_301);
    fifo_csv_dumper_302 = new("./depth302.csv");
    cstatus_csv_dumper_302 = new("./chan_status302.csv");
    fifo_monitor_302 = new(fifo_csv_dumper_302,fifo_intf_302,cstatus_csv_dumper_302);
    fifo_csv_dumper_303 = new("./depth303.csv");
    cstatus_csv_dumper_303 = new("./chan_status303.csv");
    fifo_monitor_303 = new(fifo_csv_dumper_303,fifo_intf_303,cstatus_csv_dumper_303);
    fifo_csv_dumper_304 = new("./depth304.csv");
    cstatus_csv_dumper_304 = new("./chan_status304.csv");
    fifo_monitor_304 = new(fifo_csv_dumper_304,fifo_intf_304,cstatus_csv_dumper_304);
    fifo_csv_dumper_305 = new("./depth305.csv");
    cstatus_csv_dumper_305 = new("./chan_status305.csv");
    fifo_monitor_305 = new(fifo_csv_dumper_305,fifo_intf_305,cstatus_csv_dumper_305);
    fifo_csv_dumper_306 = new("./depth306.csv");
    cstatus_csv_dumper_306 = new("./chan_status306.csv");
    fifo_monitor_306 = new(fifo_csv_dumper_306,fifo_intf_306,cstatus_csv_dumper_306);
    fifo_csv_dumper_307 = new("./depth307.csv");
    cstatus_csv_dumper_307 = new("./chan_status307.csv");
    fifo_monitor_307 = new(fifo_csv_dumper_307,fifo_intf_307,cstatus_csv_dumper_307);
    fifo_csv_dumper_308 = new("./depth308.csv");
    cstatus_csv_dumper_308 = new("./chan_status308.csv");
    fifo_monitor_308 = new(fifo_csv_dumper_308,fifo_intf_308,cstatus_csv_dumper_308);
    fifo_csv_dumper_309 = new("./depth309.csv");
    cstatus_csv_dumper_309 = new("./chan_status309.csv");
    fifo_monitor_309 = new(fifo_csv_dumper_309,fifo_intf_309,cstatus_csv_dumper_309);
    fifo_csv_dumper_310 = new("./depth310.csv");
    cstatus_csv_dumper_310 = new("./chan_status310.csv");
    fifo_monitor_310 = new(fifo_csv_dumper_310,fifo_intf_310,cstatus_csv_dumper_310);
    fifo_csv_dumper_311 = new("./depth311.csv");
    cstatus_csv_dumper_311 = new("./chan_status311.csv");
    fifo_monitor_311 = new(fifo_csv_dumper_311,fifo_intf_311,cstatus_csv_dumper_311);
    fifo_csv_dumper_312 = new("./depth312.csv");
    cstatus_csv_dumper_312 = new("./chan_status312.csv");
    fifo_monitor_312 = new(fifo_csv_dumper_312,fifo_intf_312,cstatus_csv_dumper_312);
    fifo_csv_dumper_313 = new("./depth313.csv");
    cstatus_csv_dumper_313 = new("./chan_status313.csv");
    fifo_monitor_313 = new(fifo_csv_dumper_313,fifo_intf_313,cstatus_csv_dumper_313);
    fifo_csv_dumper_314 = new("./depth314.csv");
    cstatus_csv_dumper_314 = new("./chan_status314.csv");
    fifo_monitor_314 = new(fifo_csv_dumper_314,fifo_intf_314,cstatus_csv_dumper_314);
    fifo_csv_dumper_315 = new("./depth315.csv");
    cstatus_csv_dumper_315 = new("./chan_status315.csv");
    fifo_monitor_315 = new(fifo_csv_dumper_315,fifo_intf_315,cstatus_csv_dumper_315);
    fifo_csv_dumper_316 = new("./depth316.csv");
    cstatus_csv_dumper_316 = new("./chan_status316.csv");
    fifo_monitor_316 = new(fifo_csv_dumper_316,fifo_intf_316,cstatus_csv_dumper_316);
    fifo_csv_dumper_317 = new("./depth317.csv");
    cstatus_csv_dumper_317 = new("./chan_status317.csv");
    fifo_monitor_317 = new(fifo_csv_dumper_317,fifo_intf_317,cstatus_csv_dumper_317);
    fifo_csv_dumper_318 = new("./depth318.csv");
    cstatus_csv_dumper_318 = new("./chan_status318.csv");
    fifo_monitor_318 = new(fifo_csv_dumper_318,fifo_intf_318,cstatus_csv_dumper_318);
    fifo_csv_dumper_319 = new("./depth319.csv");
    cstatus_csv_dumper_319 = new("./chan_status319.csv");
    fifo_monitor_319 = new(fifo_csv_dumper_319,fifo_intf_319,cstatus_csv_dumper_319);
    fifo_csv_dumper_320 = new("./depth320.csv");
    cstatus_csv_dumper_320 = new("./chan_status320.csv");
    fifo_monitor_320 = new(fifo_csv_dumper_320,fifo_intf_320,cstatus_csv_dumper_320);
    fifo_csv_dumper_321 = new("./depth321.csv");
    cstatus_csv_dumper_321 = new("./chan_status321.csv");
    fifo_monitor_321 = new(fifo_csv_dumper_321,fifo_intf_321,cstatus_csv_dumper_321);
    fifo_csv_dumper_322 = new("./depth322.csv");
    cstatus_csv_dumper_322 = new("./chan_status322.csv");
    fifo_monitor_322 = new(fifo_csv_dumper_322,fifo_intf_322,cstatus_csv_dumper_322);
    fifo_csv_dumper_323 = new("./depth323.csv");
    cstatus_csv_dumper_323 = new("./chan_status323.csv");
    fifo_monitor_323 = new(fifo_csv_dumper_323,fifo_intf_323,cstatus_csv_dumper_323);
    fifo_csv_dumper_324 = new("./depth324.csv");
    cstatus_csv_dumper_324 = new("./chan_status324.csv");
    fifo_monitor_324 = new(fifo_csv_dumper_324,fifo_intf_324,cstatus_csv_dumper_324);
    fifo_csv_dumper_325 = new("./depth325.csv");
    cstatus_csv_dumper_325 = new("./chan_status325.csv");
    fifo_monitor_325 = new(fifo_csv_dumper_325,fifo_intf_325,cstatus_csv_dumper_325);
    fifo_csv_dumper_326 = new("./depth326.csv");
    cstatus_csv_dumper_326 = new("./chan_status326.csv");
    fifo_monitor_326 = new(fifo_csv_dumper_326,fifo_intf_326,cstatus_csv_dumper_326);
    fifo_csv_dumper_327 = new("./depth327.csv");
    cstatus_csv_dumper_327 = new("./chan_status327.csv");
    fifo_monitor_327 = new(fifo_csv_dumper_327,fifo_intf_327,cstatus_csv_dumper_327);
    fifo_csv_dumper_328 = new("./depth328.csv");
    cstatus_csv_dumper_328 = new("./chan_status328.csv");
    fifo_monitor_328 = new(fifo_csv_dumper_328,fifo_intf_328,cstatus_csv_dumper_328);
    fifo_csv_dumper_329 = new("./depth329.csv");
    cstatus_csv_dumper_329 = new("./chan_status329.csv");
    fifo_monitor_329 = new(fifo_csv_dumper_329,fifo_intf_329,cstatus_csv_dumper_329);
    fifo_csv_dumper_330 = new("./depth330.csv");
    cstatus_csv_dumper_330 = new("./chan_status330.csv");
    fifo_monitor_330 = new(fifo_csv_dumper_330,fifo_intf_330,cstatus_csv_dumper_330);
    fifo_csv_dumper_331 = new("./depth331.csv");
    cstatus_csv_dumper_331 = new("./chan_status331.csv");
    fifo_monitor_331 = new(fifo_csv_dumper_331,fifo_intf_331,cstatus_csv_dumper_331);
    fifo_csv_dumper_332 = new("./depth332.csv");
    cstatus_csv_dumper_332 = new("./chan_status332.csv");
    fifo_monitor_332 = new(fifo_csv_dumper_332,fifo_intf_332,cstatus_csv_dumper_332);
    fifo_csv_dumper_333 = new("./depth333.csv");
    cstatus_csv_dumper_333 = new("./chan_status333.csv");
    fifo_monitor_333 = new(fifo_csv_dumper_333,fifo_intf_333,cstatus_csv_dumper_333);
    fifo_csv_dumper_334 = new("./depth334.csv");
    cstatus_csv_dumper_334 = new("./chan_status334.csv");
    fifo_monitor_334 = new(fifo_csv_dumper_334,fifo_intf_334,cstatus_csv_dumper_334);
    fifo_csv_dumper_335 = new("./depth335.csv");
    cstatus_csv_dumper_335 = new("./chan_status335.csv");
    fifo_monitor_335 = new(fifo_csv_dumper_335,fifo_intf_335,cstatus_csv_dumper_335);
    fifo_csv_dumper_336 = new("./depth336.csv");
    cstatus_csv_dumper_336 = new("./chan_status336.csv");
    fifo_monitor_336 = new(fifo_csv_dumper_336,fifo_intf_336,cstatus_csv_dumper_336);
    fifo_csv_dumper_337 = new("./depth337.csv");
    cstatus_csv_dumper_337 = new("./chan_status337.csv");
    fifo_monitor_337 = new(fifo_csv_dumper_337,fifo_intf_337,cstatus_csv_dumper_337);
    fifo_csv_dumper_338 = new("./depth338.csv");
    cstatus_csv_dumper_338 = new("./chan_status338.csv");
    fifo_monitor_338 = new(fifo_csv_dumper_338,fifo_intf_338,cstatus_csv_dumper_338);
    fifo_csv_dumper_339 = new("./depth339.csv");
    cstatus_csv_dumper_339 = new("./chan_status339.csv");
    fifo_monitor_339 = new(fifo_csv_dumper_339,fifo_intf_339,cstatus_csv_dumper_339);
    fifo_csv_dumper_340 = new("./depth340.csv");
    cstatus_csv_dumper_340 = new("./chan_status340.csv");
    fifo_monitor_340 = new(fifo_csv_dumper_340,fifo_intf_340,cstatus_csv_dumper_340);
    fifo_csv_dumper_341 = new("./depth341.csv");
    cstatus_csv_dumper_341 = new("./chan_status341.csv");
    fifo_monitor_341 = new(fifo_csv_dumper_341,fifo_intf_341,cstatus_csv_dumper_341);
    fifo_csv_dumper_342 = new("./depth342.csv");
    cstatus_csv_dumper_342 = new("./chan_status342.csv");
    fifo_monitor_342 = new(fifo_csv_dumper_342,fifo_intf_342,cstatus_csv_dumper_342);
    fifo_csv_dumper_343 = new("./depth343.csv");
    cstatus_csv_dumper_343 = new("./chan_status343.csv");
    fifo_monitor_343 = new(fifo_csv_dumper_343,fifo_intf_343,cstatus_csv_dumper_343);
    fifo_csv_dumper_344 = new("./depth344.csv");
    cstatus_csv_dumper_344 = new("./chan_status344.csv");
    fifo_monitor_344 = new(fifo_csv_dumper_344,fifo_intf_344,cstatus_csv_dumper_344);
    fifo_csv_dumper_345 = new("./depth345.csv");
    cstatus_csv_dumper_345 = new("./chan_status345.csv");
    fifo_monitor_345 = new(fifo_csv_dumper_345,fifo_intf_345,cstatus_csv_dumper_345);
    fifo_csv_dumper_346 = new("./depth346.csv");
    cstatus_csv_dumper_346 = new("./chan_status346.csv");
    fifo_monitor_346 = new(fifo_csv_dumper_346,fifo_intf_346,cstatus_csv_dumper_346);
    fifo_csv_dumper_347 = new("./depth347.csv");
    cstatus_csv_dumper_347 = new("./chan_status347.csv");
    fifo_monitor_347 = new(fifo_csv_dumper_347,fifo_intf_347,cstatus_csv_dumper_347);
    fifo_csv_dumper_348 = new("./depth348.csv");
    cstatus_csv_dumper_348 = new("./chan_status348.csv");
    fifo_monitor_348 = new(fifo_csv_dumper_348,fifo_intf_348,cstatus_csv_dumper_348);
    fifo_csv_dumper_349 = new("./depth349.csv");
    cstatus_csv_dumper_349 = new("./chan_status349.csv");
    fifo_monitor_349 = new(fifo_csv_dumper_349,fifo_intf_349,cstatus_csv_dumper_349);
    fifo_csv_dumper_350 = new("./depth350.csv");
    cstatus_csv_dumper_350 = new("./chan_status350.csv");
    fifo_monitor_350 = new(fifo_csv_dumper_350,fifo_intf_350,cstatus_csv_dumper_350);
    fifo_csv_dumper_351 = new("./depth351.csv");
    cstatus_csv_dumper_351 = new("./chan_status351.csv");
    fifo_monitor_351 = new(fifo_csv_dumper_351,fifo_intf_351,cstatus_csv_dumper_351);
    fifo_csv_dumper_352 = new("./depth352.csv");
    cstatus_csv_dumper_352 = new("./chan_status352.csv");
    fifo_monitor_352 = new(fifo_csv_dumper_352,fifo_intf_352,cstatus_csv_dumper_352);
    fifo_csv_dumper_353 = new("./depth353.csv");
    cstatus_csv_dumper_353 = new("./chan_status353.csv");
    fifo_monitor_353 = new(fifo_csv_dumper_353,fifo_intf_353,cstatus_csv_dumper_353);
    fifo_csv_dumper_354 = new("./depth354.csv");
    cstatus_csv_dumper_354 = new("./chan_status354.csv");
    fifo_monitor_354 = new(fifo_csv_dumper_354,fifo_intf_354,cstatus_csv_dumper_354);
    fifo_csv_dumper_355 = new("./depth355.csv");
    cstatus_csv_dumper_355 = new("./chan_status355.csv");
    fifo_monitor_355 = new(fifo_csv_dumper_355,fifo_intf_355,cstatus_csv_dumper_355);
    fifo_csv_dumper_356 = new("./depth356.csv");
    cstatus_csv_dumper_356 = new("./chan_status356.csv");
    fifo_monitor_356 = new(fifo_csv_dumper_356,fifo_intf_356,cstatus_csv_dumper_356);
    fifo_csv_dumper_357 = new("./depth357.csv");
    cstatus_csv_dumper_357 = new("./chan_status357.csv");
    fifo_monitor_357 = new(fifo_csv_dumper_357,fifo_intf_357,cstatus_csv_dumper_357);
    fifo_csv_dumper_358 = new("./depth358.csv");
    cstatus_csv_dumper_358 = new("./chan_status358.csv");
    fifo_monitor_358 = new(fifo_csv_dumper_358,fifo_intf_358,cstatus_csv_dumper_358);
    fifo_csv_dumper_359 = new("./depth359.csv");
    cstatus_csv_dumper_359 = new("./chan_status359.csv");
    fifo_monitor_359 = new(fifo_csv_dumper_359,fifo_intf_359,cstatus_csv_dumper_359);
    fifo_csv_dumper_360 = new("./depth360.csv");
    cstatus_csv_dumper_360 = new("./chan_status360.csv");
    fifo_monitor_360 = new(fifo_csv_dumper_360,fifo_intf_360,cstatus_csv_dumper_360);
    fifo_csv_dumper_361 = new("./depth361.csv");
    cstatus_csv_dumper_361 = new("./chan_status361.csv");
    fifo_monitor_361 = new(fifo_csv_dumper_361,fifo_intf_361,cstatus_csv_dumper_361);
    fifo_csv_dumper_362 = new("./depth362.csv");
    cstatus_csv_dumper_362 = new("./chan_status362.csv");
    fifo_monitor_362 = new(fifo_csv_dumper_362,fifo_intf_362,cstatus_csv_dumper_362);
    fifo_csv_dumper_363 = new("./depth363.csv");
    cstatus_csv_dumper_363 = new("./chan_status363.csv");
    fifo_monitor_363 = new(fifo_csv_dumper_363,fifo_intf_363,cstatus_csv_dumper_363);
    fifo_csv_dumper_364 = new("./depth364.csv");
    cstatus_csv_dumper_364 = new("./chan_status364.csv");
    fifo_monitor_364 = new(fifo_csv_dumper_364,fifo_intf_364,cstatus_csv_dumper_364);
    fifo_csv_dumper_365 = new("./depth365.csv");
    cstatus_csv_dumper_365 = new("./chan_status365.csv");
    fifo_monitor_365 = new(fifo_csv_dumper_365,fifo_intf_365,cstatus_csv_dumper_365);
    fifo_csv_dumper_366 = new("./depth366.csv");
    cstatus_csv_dumper_366 = new("./chan_status366.csv");
    fifo_monitor_366 = new(fifo_csv_dumper_366,fifo_intf_366,cstatus_csv_dumper_366);
    fifo_csv_dumper_367 = new("./depth367.csv");
    cstatus_csv_dumper_367 = new("./chan_status367.csv");
    fifo_monitor_367 = new(fifo_csv_dumper_367,fifo_intf_367,cstatus_csv_dumper_367);
    fifo_csv_dumper_368 = new("./depth368.csv");
    cstatus_csv_dumper_368 = new("./chan_status368.csv");
    fifo_monitor_368 = new(fifo_csv_dumper_368,fifo_intf_368,cstatus_csv_dumper_368);
    fifo_csv_dumper_369 = new("./depth369.csv");
    cstatus_csv_dumper_369 = new("./chan_status369.csv");
    fifo_monitor_369 = new(fifo_csv_dumper_369,fifo_intf_369,cstatus_csv_dumper_369);
    fifo_csv_dumper_370 = new("./depth370.csv");
    cstatus_csv_dumper_370 = new("./chan_status370.csv");
    fifo_monitor_370 = new(fifo_csv_dumper_370,fifo_intf_370,cstatus_csv_dumper_370);
    fifo_csv_dumper_371 = new("./depth371.csv");
    cstatus_csv_dumper_371 = new("./chan_status371.csv");
    fifo_monitor_371 = new(fifo_csv_dumper_371,fifo_intf_371,cstatus_csv_dumper_371);
    fifo_csv_dumper_372 = new("./depth372.csv");
    cstatus_csv_dumper_372 = new("./chan_status372.csv");
    fifo_monitor_372 = new(fifo_csv_dumper_372,fifo_intf_372,cstatus_csv_dumper_372);
    fifo_csv_dumper_373 = new("./depth373.csv");
    cstatus_csv_dumper_373 = new("./chan_status373.csv");
    fifo_monitor_373 = new(fifo_csv_dumper_373,fifo_intf_373,cstatus_csv_dumper_373);
    fifo_csv_dumper_374 = new("./depth374.csv");
    cstatus_csv_dumper_374 = new("./chan_status374.csv");
    fifo_monitor_374 = new(fifo_csv_dumper_374,fifo_intf_374,cstatus_csv_dumper_374);
    fifo_csv_dumper_375 = new("./depth375.csv");
    cstatus_csv_dumper_375 = new("./chan_status375.csv");
    fifo_monitor_375 = new(fifo_csv_dumper_375,fifo_intf_375,cstatus_csv_dumper_375);
    fifo_csv_dumper_376 = new("./depth376.csv");
    cstatus_csv_dumper_376 = new("./chan_status376.csv");
    fifo_monitor_376 = new(fifo_csv_dumper_376,fifo_intf_376,cstatus_csv_dumper_376);
    fifo_csv_dumper_377 = new("./depth377.csv");
    cstatus_csv_dumper_377 = new("./chan_status377.csv");
    fifo_monitor_377 = new(fifo_csv_dumper_377,fifo_intf_377,cstatus_csv_dumper_377);
    fifo_csv_dumper_378 = new("./depth378.csv");
    cstatus_csv_dumper_378 = new("./chan_status378.csv");
    fifo_monitor_378 = new(fifo_csv_dumper_378,fifo_intf_378,cstatus_csv_dumper_378);
    fifo_csv_dumper_379 = new("./depth379.csv");
    cstatus_csv_dumper_379 = new("./chan_status379.csv");
    fifo_monitor_379 = new(fifo_csv_dumper_379,fifo_intf_379,cstatus_csv_dumper_379);
    fifo_csv_dumper_380 = new("./depth380.csv");
    cstatus_csv_dumper_380 = new("./chan_status380.csv");
    fifo_monitor_380 = new(fifo_csv_dumper_380,fifo_intf_380,cstatus_csv_dumper_380);
    fifo_csv_dumper_381 = new("./depth381.csv");
    cstatus_csv_dumper_381 = new("./chan_status381.csv");
    fifo_monitor_381 = new(fifo_csv_dumper_381,fifo_intf_381,cstatus_csv_dumper_381);
    fifo_csv_dumper_382 = new("./depth382.csv");
    cstatus_csv_dumper_382 = new("./chan_status382.csv");
    fifo_monitor_382 = new(fifo_csv_dumper_382,fifo_intf_382,cstatus_csv_dumper_382);
    fifo_csv_dumper_383 = new("./depth383.csv");
    cstatus_csv_dumper_383 = new("./chan_status383.csv");
    fifo_monitor_383 = new(fifo_csv_dumper_383,fifo_intf_383,cstatus_csv_dumper_383);
    fifo_csv_dumper_384 = new("./depth384.csv");
    cstatus_csv_dumper_384 = new("./chan_status384.csv");
    fifo_monitor_384 = new(fifo_csv_dumper_384,fifo_intf_384,cstatus_csv_dumper_384);
    fifo_csv_dumper_385 = new("./depth385.csv");
    cstatus_csv_dumper_385 = new("./chan_status385.csv");
    fifo_monitor_385 = new(fifo_csv_dumper_385,fifo_intf_385,cstatus_csv_dumper_385);
    fifo_csv_dumper_386 = new("./depth386.csv");
    cstatus_csv_dumper_386 = new("./chan_status386.csv");
    fifo_monitor_386 = new(fifo_csv_dumper_386,fifo_intf_386,cstatus_csv_dumper_386);
    fifo_csv_dumper_387 = new("./depth387.csv");
    cstatus_csv_dumper_387 = new("./chan_status387.csv");
    fifo_monitor_387 = new(fifo_csv_dumper_387,fifo_intf_387,cstatus_csv_dumper_387);
    fifo_csv_dumper_388 = new("./depth388.csv");
    cstatus_csv_dumper_388 = new("./chan_status388.csv");
    fifo_monitor_388 = new(fifo_csv_dumper_388,fifo_intf_388,cstatus_csv_dumper_388);
    fifo_csv_dumper_389 = new("./depth389.csv");
    cstatus_csv_dumper_389 = new("./chan_status389.csv");
    fifo_monitor_389 = new(fifo_csv_dumper_389,fifo_intf_389,cstatus_csv_dumper_389);
    fifo_csv_dumper_390 = new("./depth390.csv");
    cstatus_csv_dumper_390 = new("./chan_status390.csv");
    fifo_monitor_390 = new(fifo_csv_dumper_390,fifo_intf_390,cstatus_csv_dumper_390);
    fifo_csv_dumper_391 = new("./depth391.csv");
    cstatus_csv_dumper_391 = new("./chan_status391.csv");
    fifo_monitor_391 = new(fifo_csv_dumper_391,fifo_intf_391,cstatus_csv_dumper_391);
    fifo_csv_dumper_392 = new("./depth392.csv");
    cstatus_csv_dumper_392 = new("./chan_status392.csv");
    fifo_monitor_392 = new(fifo_csv_dumper_392,fifo_intf_392,cstatus_csv_dumper_392);
    fifo_csv_dumper_393 = new("./depth393.csv");
    cstatus_csv_dumper_393 = new("./chan_status393.csv");
    fifo_monitor_393 = new(fifo_csv_dumper_393,fifo_intf_393,cstatus_csv_dumper_393);
    fifo_csv_dumper_394 = new("./depth394.csv");
    cstatus_csv_dumper_394 = new("./chan_status394.csv");
    fifo_monitor_394 = new(fifo_csv_dumper_394,fifo_intf_394,cstatus_csv_dumper_394);
    fifo_csv_dumper_395 = new("./depth395.csv");
    cstatus_csv_dumper_395 = new("./chan_status395.csv");
    fifo_monitor_395 = new(fifo_csv_dumper_395,fifo_intf_395,cstatus_csv_dumper_395);
    fifo_csv_dumper_396 = new("./depth396.csv");
    cstatus_csv_dumper_396 = new("./chan_status396.csv");
    fifo_monitor_396 = new(fifo_csv_dumper_396,fifo_intf_396,cstatus_csv_dumper_396);
    fifo_csv_dumper_397 = new("./depth397.csv");
    cstatus_csv_dumper_397 = new("./chan_status397.csv");
    fifo_monitor_397 = new(fifo_csv_dumper_397,fifo_intf_397,cstatus_csv_dumper_397);
    fifo_csv_dumper_398 = new("./depth398.csv");
    cstatus_csv_dumper_398 = new("./chan_status398.csv");
    fifo_monitor_398 = new(fifo_csv_dumper_398,fifo_intf_398,cstatus_csv_dumper_398);
    fifo_csv_dumper_399 = new("./depth399.csv");
    cstatus_csv_dumper_399 = new("./chan_status399.csv");
    fifo_monitor_399 = new(fifo_csv_dumper_399,fifo_intf_399,cstatus_csv_dumper_399);
    fifo_csv_dumper_400 = new("./depth400.csv");
    cstatus_csv_dumper_400 = new("./chan_status400.csv");
    fifo_monitor_400 = new(fifo_csv_dumper_400,fifo_intf_400,cstatus_csv_dumper_400);
    fifo_csv_dumper_401 = new("./depth401.csv");
    cstatus_csv_dumper_401 = new("./chan_status401.csv");
    fifo_monitor_401 = new(fifo_csv_dumper_401,fifo_intf_401,cstatus_csv_dumper_401);
    fifo_csv_dumper_402 = new("./depth402.csv");
    cstatus_csv_dumper_402 = new("./chan_status402.csv");
    fifo_monitor_402 = new(fifo_csv_dumper_402,fifo_intf_402,cstatus_csv_dumper_402);
    fifo_csv_dumper_403 = new("./depth403.csv");
    cstatus_csv_dumper_403 = new("./chan_status403.csv");
    fifo_monitor_403 = new(fifo_csv_dumper_403,fifo_intf_403,cstatus_csv_dumper_403);
    fifo_csv_dumper_404 = new("./depth404.csv");
    cstatus_csv_dumper_404 = new("./chan_status404.csv");
    fifo_monitor_404 = new(fifo_csv_dumper_404,fifo_intf_404,cstatus_csv_dumper_404);
    fifo_csv_dumper_405 = new("./depth405.csv");
    cstatus_csv_dumper_405 = new("./chan_status405.csv");
    fifo_monitor_405 = new(fifo_csv_dumper_405,fifo_intf_405,cstatus_csv_dumper_405);
    fifo_csv_dumper_406 = new("./depth406.csv");
    cstatus_csv_dumper_406 = new("./chan_status406.csv");
    fifo_monitor_406 = new(fifo_csv_dumper_406,fifo_intf_406,cstatus_csv_dumper_406);
    fifo_csv_dumper_407 = new("./depth407.csv");
    cstatus_csv_dumper_407 = new("./chan_status407.csv");
    fifo_monitor_407 = new(fifo_csv_dumper_407,fifo_intf_407,cstatus_csv_dumper_407);
    fifo_csv_dumper_408 = new("./depth408.csv");
    cstatus_csv_dumper_408 = new("./chan_status408.csv");
    fifo_monitor_408 = new(fifo_csv_dumper_408,fifo_intf_408,cstatus_csv_dumper_408);
    fifo_csv_dumper_409 = new("./depth409.csv");
    cstatus_csv_dumper_409 = new("./chan_status409.csv");
    fifo_monitor_409 = new(fifo_csv_dumper_409,fifo_intf_409,cstatus_csv_dumper_409);
    fifo_csv_dumper_410 = new("./depth410.csv");
    cstatus_csv_dumper_410 = new("./chan_status410.csv");
    fifo_monitor_410 = new(fifo_csv_dumper_410,fifo_intf_410,cstatus_csv_dumper_410);
    fifo_csv_dumper_411 = new("./depth411.csv");
    cstatus_csv_dumper_411 = new("./chan_status411.csv");
    fifo_monitor_411 = new(fifo_csv_dumper_411,fifo_intf_411,cstatus_csv_dumper_411);
    fifo_csv_dumper_412 = new("./depth412.csv");
    cstatus_csv_dumper_412 = new("./chan_status412.csv");
    fifo_monitor_412 = new(fifo_csv_dumper_412,fifo_intf_412,cstatus_csv_dumper_412);
    fifo_csv_dumper_413 = new("./depth413.csv");
    cstatus_csv_dumper_413 = new("./chan_status413.csv");
    fifo_monitor_413 = new(fifo_csv_dumper_413,fifo_intf_413,cstatus_csv_dumper_413);
    fifo_csv_dumper_414 = new("./depth414.csv");
    cstatus_csv_dumper_414 = new("./chan_status414.csv");
    fifo_monitor_414 = new(fifo_csv_dumper_414,fifo_intf_414,cstatus_csv_dumper_414);
    fifo_csv_dumper_415 = new("./depth415.csv");
    cstatus_csv_dumper_415 = new("./chan_status415.csv");
    fifo_monitor_415 = new(fifo_csv_dumper_415,fifo_intf_415,cstatus_csv_dumper_415);
    fifo_csv_dumper_416 = new("./depth416.csv");
    cstatus_csv_dumper_416 = new("./chan_status416.csv");
    fifo_monitor_416 = new(fifo_csv_dumper_416,fifo_intf_416,cstatus_csv_dumper_416);
    fifo_csv_dumper_417 = new("./depth417.csv");
    cstatus_csv_dumper_417 = new("./chan_status417.csv");
    fifo_monitor_417 = new(fifo_csv_dumper_417,fifo_intf_417,cstatus_csv_dumper_417);
    fifo_csv_dumper_418 = new("./depth418.csv");
    cstatus_csv_dumper_418 = new("./chan_status418.csv");
    fifo_monitor_418 = new(fifo_csv_dumper_418,fifo_intf_418,cstatus_csv_dumper_418);
    fifo_csv_dumper_419 = new("./depth419.csv");
    cstatus_csv_dumper_419 = new("./chan_status419.csv");
    fifo_monitor_419 = new(fifo_csv_dumper_419,fifo_intf_419,cstatus_csv_dumper_419);
    fifo_csv_dumper_420 = new("./depth420.csv");
    cstatus_csv_dumper_420 = new("./chan_status420.csv");
    fifo_monitor_420 = new(fifo_csv_dumper_420,fifo_intf_420,cstatus_csv_dumper_420);
    fifo_csv_dumper_421 = new("./depth421.csv");
    cstatus_csv_dumper_421 = new("./chan_status421.csv");
    fifo_monitor_421 = new(fifo_csv_dumper_421,fifo_intf_421,cstatus_csv_dumper_421);
    fifo_csv_dumper_422 = new("./depth422.csv");
    cstatus_csv_dumper_422 = new("./chan_status422.csv");
    fifo_monitor_422 = new(fifo_csv_dumper_422,fifo_intf_422,cstatus_csv_dumper_422);
    fifo_csv_dumper_423 = new("./depth423.csv");
    cstatus_csv_dumper_423 = new("./chan_status423.csv");
    fifo_monitor_423 = new(fifo_csv_dumper_423,fifo_intf_423,cstatus_csv_dumper_423);
    fifo_csv_dumper_424 = new("./depth424.csv");
    cstatus_csv_dumper_424 = new("./chan_status424.csv");
    fifo_monitor_424 = new(fifo_csv_dumper_424,fifo_intf_424,cstatus_csv_dumper_424);
    fifo_csv_dumper_425 = new("./depth425.csv");
    cstatus_csv_dumper_425 = new("./chan_status425.csv");
    fifo_monitor_425 = new(fifo_csv_dumper_425,fifo_intf_425,cstatus_csv_dumper_425);
    fifo_csv_dumper_426 = new("./depth426.csv");
    cstatus_csv_dumper_426 = new("./chan_status426.csv");
    fifo_monitor_426 = new(fifo_csv_dumper_426,fifo_intf_426,cstatus_csv_dumper_426);
    fifo_csv_dumper_427 = new("./depth427.csv");
    cstatus_csv_dumper_427 = new("./chan_status427.csv");
    fifo_monitor_427 = new(fifo_csv_dumper_427,fifo_intf_427,cstatus_csv_dumper_427);
    fifo_csv_dumper_428 = new("./depth428.csv");
    cstatus_csv_dumper_428 = new("./chan_status428.csv");
    fifo_monitor_428 = new(fifo_csv_dumper_428,fifo_intf_428,cstatus_csv_dumper_428);
    fifo_csv_dumper_429 = new("./depth429.csv");
    cstatus_csv_dumper_429 = new("./chan_status429.csv");
    fifo_monitor_429 = new(fifo_csv_dumper_429,fifo_intf_429,cstatus_csv_dumper_429);
    fifo_csv_dumper_430 = new("./depth430.csv");
    cstatus_csv_dumper_430 = new("./chan_status430.csv");
    fifo_monitor_430 = new(fifo_csv_dumper_430,fifo_intf_430,cstatus_csv_dumper_430);
    fifo_csv_dumper_431 = new("./depth431.csv");
    cstatus_csv_dumper_431 = new("./chan_status431.csv");
    fifo_monitor_431 = new(fifo_csv_dumper_431,fifo_intf_431,cstatus_csv_dumper_431);
    fifo_csv_dumper_432 = new("./depth432.csv");
    cstatus_csv_dumper_432 = new("./chan_status432.csv");
    fifo_monitor_432 = new(fifo_csv_dumper_432,fifo_intf_432,cstatus_csv_dumper_432);
    fifo_csv_dumper_433 = new("./depth433.csv");
    cstatus_csv_dumper_433 = new("./chan_status433.csv");
    fifo_monitor_433 = new(fifo_csv_dumper_433,fifo_intf_433,cstatus_csv_dumper_433);
    fifo_csv_dumper_434 = new("./depth434.csv");
    cstatus_csv_dumper_434 = new("./chan_status434.csv");
    fifo_monitor_434 = new(fifo_csv_dumper_434,fifo_intf_434,cstatus_csv_dumper_434);
    fifo_csv_dumper_435 = new("./depth435.csv");
    cstatus_csv_dumper_435 = new("./chan_status435.csv");
    fifo_monitor_435 = new(fifo_csv_dumper_435,fifo_intf_435,cstatus_csv_dumper_435);
    fifo_csv_dumper_436 = new("./depth436.csv");
    cstatus_csv_dumper_436 = new("./chan_status436.csv");
    fifo_monitor_436 = new(fifo_csv_dumper_436,fifo_intf_436,cstatus_csv_dumper_436);
    fifo_csv_dumper_437 = new("./depth437.csv");
    cstatus_csv_dumper_437 = new("./chan_status437.csv");
    fifo_monitor_437 = new(fifo_csv_dumper_437,fifo_intf_437,cstatus_csv_dumper_437);
    fifo_csv_dumper_438 = new("./depth438.csv");
    cstatus_csv_dumper_438 = new("./chan_status438.csv");
    fifo_monitor_438 = new(fifo_csv_dumper_438,fifo_intf_438,cstatus_csv_dumper_438);
    fifo_csv_dumper_439 = new("./depth439.csv");
    cstatus_csv_dumper_439 = new("./chan_status439.csv");
    fifo_monitor_439 = new(fifo_csv_dumper_439,fifo_intf_439,cstatus_csv_dumper_439);
    fifo_csv_dumper_440 = new("./depth440.csv");
    cstatus_csv_dumper_440 = new("./chan_status440.csv");
    fifo_monitor_440 = new(fifo_csv_dumper_440,fifo_intf_440,cstatus_csv_dumper_440);
    fifo_csv_dumper_441 = new("./depth441.csv");
    cstatus_csv_dumper_441 = new("./chan_status441.csv");
    fifo_monitor_441 = new(fifo_csv_dumper_441,fifo_intf_441,cstatus_csv_dumper_441);
    fifo_csv_dumper_442 = new("./depth442.csv");
    cstatus_csv_dumper_442 = new("./chan_status442.csv");
    fifo_monitor_442 = new(fifo_csv_dumper_442,fifo_intf_442,cstatus_csv_dumper_442);
    fifo_csv_dumper_443 = new("./depth443.csv");
    cstatus_csv_dumper_443 = new("./chan_status443.csv");
    fifo_monitor_443 = new(fifo_csv_dumper_443,fifo_intf_443,cstatus_csv_dumper_443);
    fifo_csv_dumper_444 = new("./depth444.csv");
    cstatus_csv_dumper_444 = new("./chan_status444.csv");
    fifo_monitor_444 = new(fifo_csv_dumper_444,fifo_intf_444,cstatus_csv_dumper_444);
    fifo_csv_dumper_445 = new("./depth445.csv");
    cstatus_csv_dumper_445 = new("./chan_status445.csv");
    fifo_monitor_445 = new(fifo_csv_dumper_445,fifo_intf_445,cstatus_csv_dumper_445);
    fifo_csv_dumper_446 = new("./depth446.csv");
    cstatus_csv_dumper_446 = new("./chan_status446.csv");
    fifo_monitor_446 = new(fifo_csv_dumper_446,fifo_intf_446,cstatus_csv_dumper_446);
    fifo_csv_dumper_447 = new("./depth447.csv");
    cstatus_csv_dumper_447 = new("./chan_status447.csv");
    fifo_monitor_447 = new(fifo_csv_dumper_447,fifo_intf_447,cstatus_csv_dumper_447);
    fifo_csv_dumper_448 = new("./depth448.csv");
    cstatus_csv_dumper_448 = new("./chan_status448.csv");
    fifo_monitor_448 = new(fifo_csv_dumper_448,fifo_intf_448,cstatus_csv_dumper_448);
    fifo_csv_dumper_449 = new("./depth449.csv");
    cstatus_csv_dumper_449 = new("./chan_status449.csv");
    fifo_monitor_449 = new(fifo_csv_dumper_449,fifo_intf_449,cstatus_csv_dumper_449);
    fifo_csv_dumper_450 = new("./depth450.csv");
    cstatus_csv_dumper_450 = new("./chan_status450.csv");
    fifo_monitor_450 = new(fifo_csv_dumper_450,fifo_intf_450,cstatus_csv_dumper_450);
    fifo_csv_dumper_451 = new("./depth451.csv");
    cstatus_csv_dumper_451 = new("./chan_status451.csv");
    fifo_monitor_451 = new(fifo_csv_dumper_451,fifo_intf_451,cstatus_csv_dumper_451);
    fifo_csv_dumper_452 = new("./depth452.csv");
    cstatus_csv_dumper_452 = new("./chan_status452.csv");
    fifo_monitor_452 = new(fifo_csv_dumper_452,fifo_intf_452,cstatus_csv_dumper_452);
    fifo_csv_dumper_453 = new("./depth453.csv");
    cstatus_csv_dumper_453 = new("./chan_status453.csv");
    fifo_monitor_453 = new(fifo_csv_dumper_453,fifo_intf_453,cstatus_csv_dumper_453);
    fifo_csv_dumper_454 = new("./depth454.csv");
    cstatus_csv_dumper_454 = new("./chan_status454.csv");
    fifo_monitor_454 = new(fifo_csv_dumper_454,fifo_intf_454,cstatus_csv_dumper_454);
    fifo_csv_dumper_455 = new("./depth455.csv");
    cstatus_csv_dumper_455 = new("./chan_status455.csv");
    fifo_monitor_455 = new(fifo_csv_dumper_455,fifo_intf_455,cstatus_csv_dumper_455);
    fifo_csv_dumper_456 = new("./depth456.csv");
    cstatus_csv_dumper_456 = new("./chan_status456.csv");
    fifo_monitor_456 = new(fifo_csv_dumper_456,fifo_intf_456,cstatus_csv_dumper_456);
    fifo_csv_dumper_457 = new("./depth457.csv");
    cstatus_csv_dumper_457 = new("./chan_status457.csv");
    fifo_monitor_457 = new(fifo_csv_dumper_457,fifo_intf_457,cstatus_csv_dumper_457);
    fifo_csv_dumper_458 = new("./depth458.csv");
    cstatus_csv_dumper_458 = new("./chan_status458.csv");
    fifo_monitor_458 = new(fifo_csv_dumper_458,fifo_intf_458,cstatus_csv_dumper_458);
    fifo_csv_dumper_459 = new("./depth459.csv");
    cstatus_csv_dumper_459 = new("./chan_status459.csv");
    fifo_monitor_459 = new(fifo_csv_dumper_459,fifo_intf_459,cstatus_csv_dumper_459);
    fifo_csv_dumper_460 = new("./depth460.csv");
    cstatus_csv_dumper_460 = new("./chan_status460.csv");
    fifo_monitor_460 = new(fifo_csv_dumper_460,fifo_intf_460,cstatus_csv_dumper_460);
    fifo_csv_dumper_461 = new("./depth461.csv");
    cstatus_csv_dumper_461 = new("./chan_status461.csv");
    fifo_monitor_461 = new(fifo_csv_dumper_461,fifo_intf_461,cstatus_csv_dumper_461);
    fifo_csv_dumper_462 = new("./depth462.csv");
    cstatus_csv_dumper_462 = new("./chan_status462.csv");
    fifo_monitor_462 = new(fifo_csv_dumper_462,fifo_intf_462,cstatus_csv_dumper_462);
    fifo_csv_dumper_463 = new("./depth463.csv");
    cstatus_csv_dumper_463 = new("./chan_status463.csv");
    fifo_monitor_463 = new(fifo_csv_dumper_463,fifo_intf_463,cstatus_csv_dumper_463);
    fifo_csv_dumper_464 = new("./depth464.csv");
    cstatus_csv_dumper_464 = new("./chan_status464.csv");
    fifo_monitor_464 = new(fifo_csv_dumper_464,fifo_intf_464,cstatus_csv_dumper_464);
    fifo_csv_dumper_465 = new("./depth465.csv");
    cstatus_csv_dumper_465 = new("./chan_status465.csv");
    fifo_monitor_465 = new(fifo_csv_dumper_465,fifo_intf_465,cstatus_csv_dumper_465);
    fifo_csv_dumper_466 = new("./depth466.csv");
    cstatus_csv_dumper_466 = new("./chan_status466.csv");
    fifo_monitor_466 = new(fifo_csv_dumper_466,fifo_intf_466,cstatus_csv_dumper_466);
    fifo_csv_dumper_467 = new("./depth467.csv");
    cstatus_csv_dumper_467 = new("./chan_status467.csv");
    fifo_monitor_467 = new(fifo_csv_dumper_467,fifo_intf_467,cstatus_csv_dumper_467);
    fifo_csv_dumper_468 = new("./depth468.csv");
    cstatus_csv_dumper_468 = new("./chan_status468.csv");
    fifo_monitor_468 = new(fifo_csv_dumper_468,fifo_intf_468,cstatus_csv_dumper_468);
    fifo_csv_dumper_469 = new("./depth469.csv");
    cstatus_csv_dumper_469 = new("./chan_status469.csv");
    fifo_monitor_469 = new(fifo_csv_dumper_469,fifo_intf_469,cstatus_csv_dumper_469);
    fifo_csv_dumper_470 = new("./depth470.csv");
    cstatus_csv_dumper_470 = new("./chan_status470.csv");
    fifo_monitor_470 = new(fifo_csv_dumper_470,fifo_intf_470,cstatus_csv_dumper_470);
    fifo_csv_dumper_471 = new("./depth471.csv");
    cstatus_csv_dumper_471 = new("./chan_status471.csv");
    fifo_monitor_471 = new(fifo_csv_dumper_471,fifo_intf_471,cstatus_csv_dumper_471);
    fifo_csv_dumper_472 = new("./depth472.csv");
    cstatus_csv_dumper_472 = new("./chan_status472.csv");
    fifo_monitor_472 = new(fifo_csv_dumper_472,fifo_intf_472,cstatus_csv_dumper_472);
    fifo_csv_dumper_473 = new("./depth473.csv");
    cstatus_csv_dumper_473 = new("./chan_status473.csv");
    fifo_monitor_473 = new(fifo_csv_dumper_473,fifo_intf_473,cstatus_csv_dumper_473);
    fifo_csv_dumper_474 = new("./depth474.csv");
    cstatus_csv_dumper_474 = new("./chan_status474.csv");
    fifo_monitor_474 = new(fifo_csv_dumper_474,fifo_intf_474,cstatus_csv_dumper_474);
    fifo_csv_dumper_475 = new("./depth475.csv");
    cstatus_csv_dumper_475 = new("./chan_status475.csv");
    fifo_monitor_475 = new(fifo_csv_dumper_475,fifo_intf_475,cstatus_csv_dumper_475);
    fifo_csv_dumper_476 = new("./depth476.csv");
    cstatus_csv_dumper_476 = new("./chan_status476.csv");
    fifo_monitor_476 = new(fifo_csv_dumper_476,fifo_intf_476,cstatus_csv_dumper_476);
    fifo_csv_dumper_477 = new("./depth477.csv");
    cstatus_csv_dumper_477 = new("./chan_status477.csv");
    fifo_monitor_477 = new(fifo_csv_dumper_477,fifo_intf_477,cstatus_csv_dumper_477);
    fifo_csv_dumper_478 = new("./depth478.csv");
    cstatus_csv_dumper_478 = new("./chan_status478.csv");
    fifo_monitor_478 = new(fifo_csv_dumper_478,fifo_intf_478,cstatus_csv_dumper_478);
    fifo_csv_dumper_479 = new("./depth479.csv");
    cstatus_csv_dumper_479 = new("./chan_status479.csv");
    fifo_monitor_479 = new(fifo_csv_dumper_479,fifo_intf_479,cstatus_csv_dumper_479);
    fifo_csv_dumper_480 = new("./depth480.csv");
    cstatus_csv_dumper_480 = new("./chan_status480.csv");
    fifo_monitor_480 = new(fifo_csv_dumper_480,fifo_intf_480,cstatus_csv_dumper_480);
    fifo_csv_dumper_481 = new("./depth481.csv");
    cstatus_csv_dumper_481 = new("./chan_status481.csv");
    fifo_monitor_481 = new(fifo_csv_dumper_481,fifo_intf_481,cstatus_csv_dumper_481);
    fifo_csv_dumper_482 = new("./depth482.csv");
    cstatus_csv_dumper_482 = new("./chan_status482.csv");
    fifo_monitor_482 = new(fifo_csv_dumper_482,fifo_intf_482,cstatus_csv_dumper_482);
    fifo_csv_dumper_483 = new("./depth483.csv");
    cstatus_csv_dumper_483 = new("./chan_status483.csv");
    fifo_monitor_483 = new(fifo_csv_dumper_483,fifo_intf_483,cstatus_csv_dumper_483);
    fifo_csv_dumper_484 = new("./depth484.csv");
    cstatus_csv_dumper_484 = new("./chan_status484.csv");
    fifo_monitor_484 = new(fifo_csv_dumper_484,fifo_intf_484,cstatus_csv_dumper_484);
    fifo_csv_dumper_485 = new("./depth485.csv");
    cstatus_csv_dumper_485 = new("./chan_status485.csv");
    fifo_monitor_485 = new(fifo_csv_dumper_485,fifo_intf_485,cstatus_csv_dumper_485);
    fifo_csv_dumper_486 = new("./depth486.csv");
    cstatus_csv_dumper_486 = new("./chan_status486.csv");
    fifo_monitor_486 = new(fifo_csv_dumper_486,fifo_intf_486,cstatus_csv_dumper_486);
    fifo_csv_dumper_487 = new("./depth487.csv");
    cstatus_csv_dumper_487 = new("./chan_status487.csv");
    fifo_monitor_487 = new(fifo_csv_dumper_487,fifo_intf_487,cstatus_csv_dumper_487);
    fifo_csv_dumper_488 = new("./depth488.csv");
    cstatus_csv_dumper_488 = new("./chan_status488.csv");
    fifo_monitor_488 = new(fifo_csv_dumper_488,fifo_intf_488,cstatus_csv_dumper_488);
    fifo_csv_dumper_489 = new("./depth489.csv");
    cstatus_csv_dumper_489 = new("./chan_status489.csv");
    fifo_monitor_489 = new(fifo_csv_dumper_489,fifo_intf_489,cstatus_csv_dumper_489);
    fifo_csv_dumper_490 = new("./depth490.csv");
    cstatus_csv_dumper_490 = new("./chan_status490.csv");
    fifo_monitor_490 = new(fifo_csv_dumper_490,fifo_intf_490,cstatus_csv_dumper_490);
    fifo_csv_dumper_491 = new("./depth491.csv");
    cstatus_csv_dumper_491 = new("./chan_status491.csv");
    fifo_monitor_491 = new(fifo_csv_dumper_491,fifo_intf_491,cstatus_csv_dumper_491);
    fifo_csv_dumper_492 = new("./depth492.csv");
    cstatus_csv_dumper_492 = new("./chan_status492.csv");
    fifo_monitor_492 = new(fifo_csv_dumper_492,fifo_intf_492,cstatus_csv_dumper_492);
    fifo_csv_dumper_493 = new("./depth493.csv");
    cstatus_csv_dumper_493 = new("./chan_status493.csv");
    fifo_monitor_493 = new(fifo_csv_dumper_493,fifo_intf_493,cstatus_csv_dumper_493);
    fifo_csv_dumper_494 = new("./depth494.csv");
    cstatus_csv_dumper_494 = new("./chan_status494.csv");
    fifo_monitor_494 = new(fifo_csv_dumper_494,fifo_intf_494,cstatus_csv_dumper_494);
    fifo_csv_dumper_495 = new("./depth495.csv");
    cstatus_csv_dumper_495 = new("./chan_status495.csv");
    fifo_monitor_495 = new(fifo_csv_dumper_495,fifo_intf_495,cstatus_csv_dumper_495);
    fifo_csv_dumper_496 = new("./depth496.csv");
    cstatus_csv_dumper_496 = new("./chan_status496.csv");
    fifo_monitor_496 = new(fifo_csv_dumper_496,fifo_intf_496,cstatus_csv_dumper_496);
    fifo_csv_dumper_497 = new("./depth497.csv");
    cstatus_csv_dumper_497 = new("./chan_status497.csv");
    fifo_monitor_497 = new(fifo_csv_dumper_497,fifo_intf_497,cstatus_csv_dumper_497);
    fifo_csv_dumper_498 = new("./depth498.csv");
    cstatus_csv_dumper_498 = new("./chan_status498.csv");
    fifo_monitor_498 = new(fifo_csv_dumper_498,fifo_intf_498,cstatus_csv_dumper_498);
    fifo_csv_dumper_499 = new("./depth499.csv");
    cstatus_csv_dumper_499 = new("./chan_status499.csv");
    fifo_monitor_499 = new(fifo_csv_dumper_499,fifo_intf_499,cstatus_csv_dumper_499);
    fifo_csv_dumper_500 = new("./depth500.csv");
    cstatus_csv_dumper_500 = new("./chan_status500.csv");
    fifo_monitor_500 = new(fifo_csv_dumper_500,fifo_intf_500,cstatus_csv_dumper_500);
    fifo_csv_dumper_501 = new("./depth501.csv");
    cstatus_csv_dumper_501 = new("./chan_status501.csv");
    fifo_monitor_501 = new(fifo_csv_dumper_501,fifo_intf_501,cstatus_csv_dumper_501);
    fifo_csv_dumper_502 = new("./depth502.csv");
    cstatus_csv_dumper_502 = new("./chan_status502.csv");
    fifo_monitor_502 = new(fifo_csv_dumper_502,fifo_intf_502,cstatus_csv_dumper_502);
    fifo_csv_dumper_503 = new("./depth503.csv");
    cstatus_csv_dumper_503 = new("./chan_status503.csv");
    fifo_monitor_503 = new(fifo_csv_dumper_503,fifo_intf_503,cstatus_csv_dumper_503);
    fifo_csv_dumper_504 = new("./depth504.csv");
    cstatus_csv_dumper_504 = new("./chan_status504.csv");
    fifo_monitor_504 = new(fifo_csv_dumper_504,fifo_intf_504,cstatus_csv_dumper_504);
    fifo_csv_dumper_505 = new("./depth505.csv");
    cstatus_csv_dumper_505 = new("./chan_status505.csv");
    fifo_monitor_505 = new(fifo_csv_dumper_505,fifo_intf_505,cstatus_csv_dumper_505);
    fifo_csv_dumper_506 = new("./depth506.csv");
    cstatus_csv_dumper_506 = new("./chan_status506.csv");
    fifo_monitor_506 = new(fifo_csv_dumper_506,fifo_intf_506,cstatus_csv_dumper_506);
    fifo_csv_dumper_507 = new("./depth507.csv");
    cstatus_csv_dumper_507 = new("./chan_status507.csv");
    fifo_monitor_507 = new(fifo_csv_dumper_507,fifo_intf_507,cstatus_csv_dumper_507);
    fifo_csv_dumper_508 = new("./depth508.csv");
    cstatus_csv_dumper_508 = new("./chan_status508.csv");
    fifo_monitor_508 = new(fifo_csv_dumper_508,fifo_intf_508,cstatus_csv_dumper_508);
    fifo_csv_dumper_509 = new("./depth509.csv");
    cstatus_csv_dumper_509 = new("./chan_status509.csv");
    fifo_monitor_509 = new(fifo_csv_dumper_509,fifo_intf_509,cstatus_csv_dumper_509);
    fifo_csv_dumper_510 = new("./depth510.csv");
    cstatus_csv_dumper_510 = new("./chan_status510.csv");
    fifo_monitor_510 = new(fifo_csv_dumper_510,fifo_intf_510,cstatus_csv_dumper_510);
    fifo_csv_dumper_511 = new("./depth511.csv");
    cstatus_csv_dumper_511 = new("./chan_status511.csv");
    fifo_monitor_511 = new(fifo_csv_dumper_511,fifo_intf_511,cstatus_csv_dumper_511);
    fifo_csv_dumper_512 = new("./depth512.csv");
    cstatus_csv_dumper_512 = new("./chan_status512.csv");
    fifo_monitor_512 = new(fifo_csv_dumper_512,fifo_intf_512,cstatus_csv_dumper_512);
    fifo_csv_dumper_513 = new("./depth513.csv");
    cstatus_csv_dumper_513 = new("./chan_status513.csv");
    fifo_monitor_513 = new(fifo_csv_dumper_513,fifo_intf_513,cstatus_csv_dumper_513);
    fifo_csv_dumper_514 = new("./depth514.csv");
    cstatus_csv_dumper_514 = new("./chan_status514.csv");
    fifo_monitor_514 = new(fifo_csv_dumper_514,fifo_intf_514,cstatus_csv_dumper_514);
    fifo_csv_dumper_515 = new("./depth515.csv");
    cstatus_csv_dumper_515 = new("./chan_status515.csv");
    fifo_monitor_515 = new(fifo_csv_dumper_515,fifo_intf_515,cstatus_csv_dumper_515);
    fifo_csv_dumper_516 = new("./depth516.csv");
    cstatus_csv_dumper_516 = new("./chan_status516.csv");
    fifo_monitor_516 = new(fifo_csv_dumper_516,fifo_intf_516,cstatus_csv_dumper_516);
    fifo_csv_dumper_517 = new("./depth517.csv");
    cstatus_csv_dumper_517 = new("./chan_status517.csv");
    fifo_monitor_517 = new(fifo_csv_dumper_517,fifo_intf_517,cstatus_csv_dumper_517);
    fifo_csv_dumper_518 = new("./depth518.csv");
    cstatus_csv_dumper_518 = new("./chan_status518.csv");
    fifo_monitor_518 = new(fifo_csv_dumper_518,fifo_intf_518,cstatus_csv_dumper_518);
    fifo_csv_dumper_519 = new("./depth519.csv");
    cstatus_csv_dumper_519 = new("./chan_status519.csv");
    fifo_monitor_519 = new(fifo_csv_dumper_519,fifo_intf_519,cstatus_csv_dumper_519);
    fifo_csv_dumper_520 = new("./depth520.csv");
    cstatus_csv_dumper_520 = new("./chan_status520.csv");
    fifo_monitor_520 = new(fifo_csv_dumper_520,fifo_intf_520,cstatus_csv_dumper_520);
    fifo_csv_dumper_521 = new("./depth521.csv");
    cstatus_csv_dumper_521 = new("./chan_status521.csv");
    fifo_monitor_521 = new(fifo_csv_dumper_521,fifo_intf_521,cstatus_csv_dumper_521);
    fifo_csv_dumper_522 = new("./depth522.csv");
    cstatus_csv_dumper_522 = new("./chan_status522.csv");
    fifo_monitor_522 = new(fifo_csv_dumper_522,fifo_intf_522,cstatus_csv_dumper_522);
    fifo_csv_dumper_523 = new("./depth523.csv");
    cstatus_csv_dumper_523 = new("./chan_status523.csv");
    fifo_monitor_523 = new(fifo_csv_dumper_523,fifo_intf_523,cstatus_csv_dumper_523);
    fifo_csv_dumper_524 = new("./depth524.csv");
    cstatus_csv_dumper_524 = new("./chan_status524.csv");
    fifo_monitor_524 = new(fifo_csv_dumper_524,fifo_intf_524,cstatus_csv_dumper_524);
    fifo_csv_dumper_525 = new("./depth525.csv");
    cstatus_csv_dumper_525 = new("./chan_status525.csv");
    fifo_monitor_525 = new(fifo_csv_dumper_525,fifo_intf_525,cstatus_csv_dumper_525);
    fifo_csv_dumper_526 = new("./depth526.csv");
    cstatus_csv_dumper_526 = new("./chan_status526.csv");
    fifo_monitor_526 = new(fifo_csv_dumper_526,fifo_intf_526,cstatus_csv_dumper_526);
    fifo_csv_dumper_527 = new("./depth527.csv");
    cstatus_csv_dumper_527 = new("./chan_status527.csv");
    fifo_monitor_527 = new(fifo_csv_dumper_527,fifo_intf_527,cstatus_csv_dumper_527);
    fifo_csv_dumper_528 = new("./depth528.csv");
    cstatus_csv_dumper_528 = new("./chan_status528.csv");
    fifo_monitor_528 = new(fifo_csv_dumper_528,fifo_intf_528,cstatus_csv_dumper_528);
    fifo_csv_dumper_529 = new("./depth529.csv");
    cstatus_csv_dumper_529 = new("./chan_status529.csv");
    fifo_monitor_529 = new(fifo_csv_dumper_529,fifo_intf_529,cstatus_csv_dumper_529);
    fifo_csv_dumper_530 = new("./depth530.csv");
    cstatus_csv_dumper_530 = new("./chan_status530.csv");
    fifo_monitor_530 = new(fifo_csv_dumper_530,fifo_intf_530,cstatus_csv_dumper_530);
    fifo_csv_dumper_531 = new("./depth531.csv");
    cstatus_csv_dumper_531 = new("./chan_status531.csv");
    fifo_monitor_531 = new(fifo_csv_dumper_531,fifo_intf_531,cstatus_csv_dumper_531);
    fifo_csv_dumper_532 = new("./depth532.csv");
    cstatus_csv_dumper_532 = new("./chan_status532.csv");
    fifo_monitor_532 = new(fifo_csv_dumper_532,fifo_intf_532,cstatus_csv_dumper_532);
    fifo_csv_dumper_533 = new("./depth533.csv");
    cstatus_csv_dumper_533 = new("./chan_status533.csv");
    fifo_monitor_533 = new(fifo_csv_dumper_533,fifo_intf_533,cstatus_csv_dumper_533);
    fifo_csv_dumper_534 = new("./depth534.csv");
    cstatus_csv_dumper_534 = new("./chan_status534.csv");
    fifo_monitor_534 = new(fifo_csv_dumper_534,fifo_intf_534,cstatus_csv_dumper_534);
    fifo_csv_dumper_535 = new("./depth535.csv");
    cstatus_csv_dumper_535 = new("./chan_status535.csv");
    fifo_monitor_535 = new(fifo_csv_dumper_535,fifo_intf_535,cstatus_csv_dumper_535);
    fifo_csv_dumper_536 = new("./depth536.csv");
    cstatus_csv_dumper_536 = new("./chan_status536.csv");
    fifo_monitor_536 = new(fifo_csv_dumper_536,fifo_intf_536,cstatus_csv_dumper_536);
    fifo_csv_dumper_537 = new("./depth537.csv");
    cstatus_csv_dumper_537 = new("./chan_status537.csv");
    fifo_monitor_537 = new(fifo_csv_dumper_537,fifo_intf_537,cstatus_csv_dumper_537);
    fifo_csv_dumper_538 = new("./depth538.csv");
    cstatus_csv_dumper_538 = new("./chan_status538.csv");
    fifo_monitor_538 = new(fifo_csv_dumper_538,fifo_intf_538,cstatus_csv_dumper_538);
    fifo_csv_dumper_539 = new("./depth539.csv");
    cstatus_csv_dumper_539 = new("./chan_status539.csv");
    fifo_monitor_539 = new(fifo_csv_dumper_539,fifo_intf_539,cstatus_csv_dumper_539);
    fifo_csv_dumper_540 = new("./depth540.csv");
    cstatus_csv_dumper_540 = new("./chan_status540.csv");
    fifo_monitor_540 = new(fifo_csv_dumper_540,fifo_intf_540,cstatus_csv_dumper_540);
    fifo_csv_dumper_541 = new("./depth541.csv");
    cstatus_csv_dumper_541 = new("./chan_status541.csv");
    fifo_monitor_541 = new(fifo_csv_dumper_541,fifo_intf_541,cstatus_csv_dumper_541);
    fifo_csv_dumper_542 = new("./depth542.csv");
    cstatus_csv_dumper_542 = new("./chan_status542.csv");
    fifo_monitor_542 = new(fifo_csv_dumper_542,fifo_intf_542,cstatus_csv_dumper_542);
    fifo_csv_dumper_543 = new("./depth543.csv");
    cstatus_csv_dumper_543 = new("./chan_status543.csv");
    fifo_monitor_543 = new(fifo_csv_dumper_543,fifo_intf_543,cstatus_csv_dumper_543);
    fifo_csv_dumper_544 = new("./depth544.csv");
    cstatus_csv_dumper_544 = new("./chan_status544.csv");
    fifo_monitor_544 = new(fifo_csv_dumper_544,fifo_intf_544,cstatus_csv_dumper_544);
    fifo_csv_dumper_545 = new("./depth545.csv");
    cstatus_csv_dumper_545 = new("./chan_status545.csv");
    fifo_monitor_545 = new(fifo_csv_dumper_545,fifo_intf_545,cstatus_csv_dumper_545);
    fifo_csv_dumper_546 = new("./depth546.csv");
    cstatus_csv_dumper_546 = new("./chan_status546.csv");
    fifo_monitor_546 = new(fifo_csv_dumper_546,fifo_intf_546,cstatus_csv_dumper_546);
    fifo_csv_dumper_547 = new("./depth547.csv");
    cstatus_csv_dumper_547 = new("./chan_status547.csv");
    fifo_monitor_547 = new(fifo_csv_dumper_547,fifo_intf_547,cstatus_csv_dumper_547);
    fifo_csv_dumper_548 = new("./depth548.csv");
    cstatus_csv_dumper_548 = new("./chan_status548.csv");
    fifo_monitor_548 = new(fifo_csv_dumper_548,fifo_intf_548,cstatus_csv_dumper_548);
    fifo_csv_dumper_549 = new("./depth549.csv");
    cstatus_csv_dumper_549 = new("./chan_status549.csv");
    fifo_monitor_549 = new(fifo_csv_dumper_549,fifo_intf_549,cstatus_csv_dumper_549);
    fifo_csv_dumper_550 = new("./depth550.csv");
    cstatus_csv_dumper_550 = new("./chan_status550.csv");
    fifo_monitor_550 = new(fifo_csv_dumper_550,fifo_intf_550,cstatus_csv_dumper_550);
    fifo_csv_dumper_551 = new("./depth551.csv");
    cstatus_csv_dumper_551 = new("./chan_status551.csv");
    fifo_monitor_551 = new(fifo_csv_dumper_551,fifo_intf_551,cstatus_csv_dumper_551);
    fifo_csv_dumper_552 = new("./depth552.csv");
    cstatus_csv_dumper_552 = new("./chan_status552.csv");
    fifo_monitor_552 = new(fifo_csv_dumper_552,fifo_intf_552,cstatus_csv_dumper_552);
    fifo_csv_dumper_553 = new("./depth553.csv");
    cstatus_csv_dumper_553 = new("./chan_status553.csv");
    fifo_monitor_553 = new(fifo_csv_dumper_553,fifo_intf_553,cstatus_csv_dumper_553);
    fifo_csv_dumper_554 = new("./depth554.csv");
    cstatus_csv_dumper_554 = new("./chan_status554.csv");
    fifo_monitor_554 = new(fifo_csv_dumper_554,fifo_intf_554,cstatus_csv_dumper_554);
    fifo_csv_dumper_555 = new("./depth555.csv");
    cstatus_csv_dumper_555 = new("./chan_status555.csv");
    fifo_monitor_555 = new(fifo_csv_dumper_555,fifo_intf_555,cstatus_csv_dumper_555);
    fifo_csv_dumper_556 = new("./depth556.csv");
    cstatus_csv_dumper_556 = new("./chan_status556.csv");
    fifo_monitor_556 = new(fifo_csv_dumper_556,fifo_intf_556,cstatus_csv_dumper_556);
    fifo_csv_dumper_557 = new("./depth557.csv");
    cstatus_csv_dumper_557 = new("./chan_status557.csv");
    fifo_monitor_557 = new(fifo_csv_dumper_557,fifo_intf_557,cstatus_csv_dumper_557);
    fifo_csv_dumper_558 = new("./depth558.csv");
    cstatus_csv_dumper_558 = new("./chan_status558.csv");
    fifo_monitor_558 = new(fifo_csv_dumper_558,fifo_intf_558,cstatus_csv_dumper_558);
    fifo_csv_dumper_559 = new("./depth559.csv");
    cstatus_csv_dumper_559 = new("./chan_status559.csv");
    fifo_monitor_559 = new(fifo_csv_dumper_559,fifo_intf_559,cstatus_csv_dumper_559);
    fifo_csv_dumper_560 = new("./depth560.csv");
    cstatus_csv_dumper_560 = new("./chan_status560.csv");
    fifo_monitor_560 = new(fifo_csv_dumper_560,fifo_intf_560,cstatus_csv_dumper_560);
    fifo_csv_dumper_561 = new("./depth561.csv");
    cstatus_csv_dumper_561 = new("./chan_status561.csv");
    fifo_monitor_561 = new(fifo_csv_dumper_561,fifo_intf_561,cstatus_csv_dumper_561);
    fifo_csv_dumper_562 = new("./depth562.csv");
    cstatus_csv_dumper_562 = new("./chan_status562.csv");
    fifo_monitor_562 = new(fifo_csv_dumper_562,fifo_intf_562,cstatus_csv_dumper_562);
    fifo_csv_dumper_563 = new("./depth563.csv");
    cstatus_csv_dumper_563 = new("./chan_status563.csv");
    fifo_monitor_563 = new(fifo_csv_dumper_563,fifo_intf_563,cstatus_csv_dumper_563);
    fifo_csv_dumper_564 = new("./depth564.csv");
    cstatus_csv_dumper_564 = new("./chan_status564.csv");
    fifo_monitor_564 = new(fifo_csv_dumper_564,fifo_intf_564,cstatus_csv_dumper_564);
    fifo_csv_dumper_565 = new("./depth565.csv");
    cstatus_csv_dumper_565 = new("./chan_status565.csv");
    fifo_monitor_565 = new(fifo_csv_dumper_565,fifo_intf_565,cstatus_csv_dumper_565);
    fifo_csv_dumper_566 = new("./depth566.csv");
    cstatus_csv_dumper_566 = new("./chan_status566.csv");
    fifo_monitor_566 = new(fifo_csv_dumper_566,fifo_intf_566,cstatus_csv_dumper_566);
    fifo_csv_dumper_567 = new("./depth567.csv");
    cstatus_csv_dumper_567 = new("./chan_status567.csv");
    fifo_monitor_567 = new(fifo_csv_dumper_567,fifo_intf_567,cstatus_csv_dumper_567);
    fifo_csv_dumper_568 = new("./depth568.csv");
    cstatus_csv_dumper_568 = new("./chan_status568.csv");
    fifo_monitor_568 = new(fifo_csv_dumper_568,fifo_intf_568,cstatus_csv_dumper_568);
    fifo_csv_dumper_569 = new("./depth569.csv");
    cstatus_csv_dumper_569 = new("./chan_status569.csv");
    fifo_monitor_569 = new(fifo_csv_dumper_569,fifo_intf_569,cstatus_csv_dumper_569);
    fifo_csv_dumper_570 = new("./depth570.csv");
    cstatus_csv_dumper_570 = new("./chan_status570.csv");
    fifo_monitor_570 = new(fifo_csv_dumper_570,fifo_intf_570,cstatus_csv_dumper_570);
    fifo_csv_dumper_571 = new("./depth571.csv");
    cstatus_csv_dumper_571 = new("./chan_status571.csv");
    fifo_monitor_571 = new(fifo_csv_dumper_571,fifo_intf_571,cstatus_csv_dumper_571);
    fifo_csv_dumper_572 = new("./depth572.csv");
    cstatus_csv_dumper_572 = new("./chan_status572.csv");
    fifo_monitor_572 = new(fifo_csv_dumper_572,fifo_intf_572,cstatus_csv_dumper_572);
    fifo_csv_dumper_573 = new("./depth573.csv");
    cstatus_csv_dumper_573 = new("./chan_status573.csv");
    fifo_monitor_573 = new(fifo_csv_dumper_573,fifo_intf_573,cstatus_csv_dumper_573);
    fifo_csv_dumper_574 = new("./depth574.csv");
    cstatus_csv_dumper_574 = new("./chan_status574.csv");
    fifo_monitor_574 = new(fifo_csv_dumper_574,fifo_intf_574,cstatus_csv_dumper_574);
    fifo_csv_dumper_575 = new("./depth575.csv");
    cstatus_csv_dumper_575 = new("./chan_status575.csv");
    fifo_monitor_575 = new(fifo_csv_dumper_575,fifo_intf_575,cstatus_csv_dumper_575);
    fifo_csv_dumper_576 = new("./depth576.csv");
    cstatus_csv_dumper_576 = new("./chan_status576.csv");
    fifo_monitor_576 = new(fifo_csv_dumper_576,fifo_intf_576,cstatus_csv_dumper_576);
    fifo_csv_dumper_577 = new("./depth577.csv");
    cstatus_csv_dumper_577 = new("./chan_status577.csv");
    fifo_monitor_577 = new(fifo_csv_dumper_577,fifo_intf_577,cstatus_csv_dumper_577);
    fifo_csv_dumper_578 = new("./depth578.csv");
    cstatus_csv_dumper_578 = new("./chan_status578.csv");
    fifo_monitor_578 = new(fifo_csv_dumper_578,fifo_intf_578,cstatus_csv_dumper_578);
    fifo_csv_dumper_579 = new("./depth579.csv");
    cstatus_csv_dumper_579 = new("./chan_status579.csv");
    fifo_monitor_579 = new(fifo_csv_dumper_579,fifo_intf_579,cstatus_csv_dumper_579);
    fifo_csv_dumper_580 = new("./depth580.csv");
    cstatus_csv_dumper_580 = new("./chan_status580.csv");
    fifo_monitor_580 = new(fifo_csv_dumper_580,fifo_intf_580,cstatus_csv_dumper_580);
    fifo_csv_dumper_581 = new("./depth581.csv");
    cstatus_csv_dumper_581 = new("./chan_status581.csv");
    fifo_monitor_581 = new(fifo_csv_dumper_581,fifo_intf_581,cstatus_csv_dumper_581);
    fifo_csv_dumper_582 = new("./depth582.csv");
    cstatus_csv_dumper_582 = new("./chan_status582.csv");
    fifo_monitor_582 = new(fifo_csv_dumper_582,fifo_intf_582,cstatus_csv_dumper_582);
    fifo_csv_dumper_583 = new("./depth583.csv");
    cstatus_csv_dumper_583 = new("./chan_status583.csv");
    fifo_monitor_583 = new(fifo_csv_dumper_583,fifo_intf_583,cstatus_csv_dumper_583);
    fifo_csv_dumper_584 = new("./depth584.csv");
    cstatus_csv_dumper_584 = new("./chan_status584.csv");
    fifo_monitor_584 = new(fifo_csv_dumper_584,fifo_intf_584,cstatus_csv_dumper_584);
    fifo_csv_dumper_585 = new("./depth585.csv");
    cstatus_csv_dumper_585 = new("./chan_status585.csv");
    fifo_monitor_585 = new(fifo_csv_dumper_585,fifo_intf_585,cstatus_csv_dumper_585);
    fifo_csv_dumper_586 = new("./depth586.csv");
    cstatus_csv_dumper_586 = new("./chan_status586.csv");
    fifo_monitor_586 = new(fifo_csv_dumper_586,fifo_intf_586,cstatus_csv_dumper_586);
    fifo_csv_dumper_587 = new("./depth587.csv");
    cstatus_csv_dumper_587 = new("./chan_status587.csv");
    fifo_monitor_587 = new(fifo_csv_dumper_587,fifo_intf_587,cstatus_csv_dumper_587);
    fifo_csv_dumper_588 = new("./depth588.csv");
    cstatus_csv_dumper_588 = new("./chan_status588.csv");
    fifo_monitor_588 = new(fifo_csv_dumper_588,fifo_intf_588,cstatus_csv_dumper_588);
    fifo_csv_dumper_589 = new("./depth589.csv");
    cstatus_csv_dumper_589 = new("./chan_status589.csv");
    fifo_monitor_589 = new(fifo_csv_dumper_589,fifo_intf_589,cstatus_csv_dumper_589);
    fifo_csv_dumper_590 = new("./depth590.csv");
    cstatus_csv_dumper_590 = new("./chan_status590.csv");
    fifo_monitor_590 = new(fifo_csv_dumper_590,fifo_intf_590,cstatus_csv_dumper_590);
    fifo_csv_dumper_591 = new("./depth591.csv");
    cstatus_csv_dumper_591 = new("./chan_status591.csv");
    fifo_monitor_591 = new(fifo_csv_dumper_591,fifo_intf_591,cstatus_csv_dumper_591);
    fifo_csv_dumper_592 = new("./depth592.csv");
    cstatus_csv_dumper_592 = new("./chan_status592.csv");
    fifo_monitor_592 = new(fifo_csv_dumper_592,fifo_intf_592,cstatus_csv_dumper_592);
    fifo_csv_dumper_593 = new("./depth593.csv");
    cstatus_csv_dumper_593 = new("./chan_status593.csv");
    fifo_monitor_593 = new(fifo_csv_dumper_593,fifo_intf_593,cstatus_csv_dumper_593);
    fifo_csv_dumper_594 = new("./depth594.csv");
    cstatus_csv_dumper_594 = new("./chan_status594.csv");
    fifo_monitor_594 = new(fifo_csv_dumper_594,fifo_intf_594,cstatus_csv_dumper_594);
    fifo_csv_dumper_595 = new("./depth595.csv");
    cstatus_csv_dumper_595 = new("./chan_status595.csv");
    fifo_monitor_595 = new(fifo_csv_dumper_595,fifo_intf_595,cstatus_csv_dumper_595);
    fifo_csv_dumper_596 = new("./depth596.csv");
    cstatus_csv_dumper_596 = new("./chan_status596.csv");
    fifo_monitor_596 = new(fifo_csv_dumper_596,fifo_intf_596,cstatus_csv_dumper_596);
    fifo_csv_dumper_597 = new("./depth597.csv");
    cstatus_csv_dumper_597 = new("./chan_status597.csv");
    fifo_monitor_597 = new(fifo_csv_dumper_597,fifo_intf_597,cstatus_csv_dumper_597);
    fifo_csv_dumper_598 = new("./depth598.csv");
    cstatus_csv_dumper_598 = new("./chan_status598.csv");
    fifo_monitor_598 = new(fifo_csv_dumper_598,fifo_intf_598,cstatus_csv_dumper_598);
    fifo_csv_dumper_599 = new("./depth599.csv");
    cstatus_csv_dumper_599 = new("./chan_status599.csv");
    fifo_monitor_599 = new(fifo_csv_dumper_599,fifo_intf_599,cstatus_csv_dumper_599);
    fifo_csv_dumper_600 = new("./depth600.csv");
    cstatus_csv_dumper_600 = new("./chan_status600.csv");
    fifo_monitor_600 = new(fifo_csv_dumper_600,fifo_intf_600,cstatus_csv_dumper_600);
    fifo_csv_dumper_601 = new("./depth601.csv");
    cstatus_csv_dumper_601 = new("./chan_status601.csv");
    fifo_monitor_601 = new(fifo_csv_dumper_601,fifo_intf_601,cstatus_csv_dumper_601);
    fifo_csv_dumper_602 = new("./depth602.csv");
    cstatus_csv_dumper_602 = new("./chan_status602.csv");
    fifo_monitor_602 = new(fifo_csv_dumper_602,fifo_intf_602,cstatus_csv_dumper_602);
    fifo_csv_dumper_603 = new("./depth603.csv");
    cstatus_csv_dumper_603 = new("./chan_status603.csv");
    fifo_monitor_603 = new(fifo_csv_dumper_603,fifo_intf_603,cstatus_csv_dumper_603);
    fifo_csv_dumper_604 = new("./depth604.csv");
    cstatus_csv_dumper_604 = new("./chan_status604.csv");
    fifo_monitor_604 = new(fifo_csv_dumper_604,fifo_intf_604,cstatus_csv_dumper_604);
    fifo_csv_dumper_605 = new("./depth605.csv");
    cstatus_csv_dumper_605 = new("./chan_status605.csv");
    fifo_monitor_605 = new(fifo_csv_dumper_605,fifo_intf_605,cstatus_csv_dumper_605);
    fifo_csv_dumper_606 = new("./depth606.csv");
    cstatus_csv_dumper_606 = new("./chan_status606.csv");
    fifo_monitor_606 = new(fifo_csv_dumper_606,fifo_intf_606,cstatus_csv_dumper_606);
    fifo_csv_dumper_607 = new("./depth607.csv");
    cstatus_csv_dumper_607 = new("./chan_status607.csv");
    fifo_monitor_607 = new(fifo_csv_dumper_607,fifo_intf_607,cstatus_csv_dumper_607);
    fifo_csv_dumper_608 = new("./depth608.csv");
    cstatus_csv_dumper_608 = new("./chan_status608.csv");
    fifo_monitor_608 = new(fifo_csv_dumper_608,fifo_intf_608,cstatus_csv_dumper_608);
    fifo_csv_dumper_609 = new("./depth609.csv");
    cstatus_csv_dumper_609 = new("./chan_status609.csv");
    fifo_monitor_609 = new(fifo_csv_dumper_609,fifo_intf_609,cstatus_csv_dumper_609);
    fifo_csv_dumper_610 = new("./depth610.csv");
    cstatus_csv_dumper_610 = new("./chan_status610.csv");
    fifo_monitor_610 = new(fifo_csv_dumper_610,fifo_intf_610,cstatus_csv_dumper_610);
    fifo_csv_dumper_611 = new("./depth611.csv");
    cstatus_csv_dumper_611 = new("./chan_status611.csv");
    fifo_monitor_611 = new(fifo_csv_dumper_611,fifo_intf_611,cstatus_csv_dumper_611);
    fifo_csv_dumper_612 = new("./depth612.csv");
    cstatus_csv_dumper_612 = new("./chan_status612.csv");
    fifo_monitor_612 = new(fifo_csv_dumper_612,fifo_intf_612,cstatus_csv_dumper_612);
    fifo_csv_dumper_613 = new("./depth613.csv");
    cstatus_csv_dumper_613 = new("./chan_status613.csv");
    fifo_monitor_613 = new(fifo_csv_dumper_613,fifo_intf_613,cstatus_csv_dumper_613);
    fifo_csv_dumper_614 = new("./depth614.csv");
    cstatus_csv_dumper_614 = new("./chan_status614.csv");
    fifo_monitor_614 = new(fifo_csv_dumper_614,fifo_intf_614,cstatus_csv_dumper_614);
    fifo_csv_dumper_615 = new("./depth615.csv");
    cstatus_csv_dumper_615 = new("./chan_status615.csv");
    fifo_monitor_615 = new(fifo_csv_dumper_615,fifo_intf_615,cstatus_csv_dumper_615);
    fifo_csv_dumper_616 = new("./depth616.csv");
    cstatus_csv_dumper_616 = new("./chan_status616.csv");
    fifo_monitor_616 = new(fifo_csv_dumper_616,fifo_intf_616,cstatus_csv_dumper_616);
    fifo_csv_dumper_617 = new("./depth617.csv");
    cstatus_csv_dumper_617 = new("./chan_status617.csv");
    fifo_monitor_617 = new(fifo_csv_dumper_617,fifo_intf_617,cstatus_csv_dumper_617);
    fifo_csv_dumper_618 = new("./depth618.csv");
    cstatus_csv_dumper_618 = new("./chan_status618.csv");
    fifo_monitor_618 = new(fifo_csv_dumper_618,fifo_intf_618,cstatus_csv_dumper_618);
    fifo_csv_dumper_619 = new("./depth619.csv");
    cstatus_csv_dumper_619 = new("./chan_status619.csv");
    fifo_monitor_619 = new(fifo_csv_dumper_619,fifo_intf_619,cstatus_csv_dumper_619);
    fifo_csv_dumper_620 = new("./depth620.csv");
    cstatus_csv_dumper_620 = new("./chan_status620.csv");
    fifo_monitor_620 = new(fifo_csv_dumper_620,fifo_intf_620,cstatus_csv_dumper_620);
    fifo_csv_dumper_621 = new("./depth621.csv");
    cstatus_csv_dumper_621 = new("./chan_status621.csv");
    fifo_monitor_621 = new(fifo_csv_dumper_621,fifo_intf_621,cstatus_csv_dumper_621);
    fifo_csv_dumper_622 = new("./depth622.csv");
    cstatus_csv_dumper_622 = new("./chan_status622.csv");
    fifo_monitor_622 = new(fifo_csv_dumper_622,fifo_intf_622,cstatus_csv_dumper_622);
    fifo_csv_dumper_623 = new("./depth623.csv");
    cstatus_csv_dumper_623 = new("./chan_status623.csv");
    fifo_monitor_623 = new(fifo_csv_dumper_623,fifo_intf_623,cstatus_csv_dumper_623);
    fifo_csv_dumper_624 = new("./depth624.csv");
    cstatus_csv_dumper_624 = new("./chan_status624.csv");
    fifo_monitor_624 = new(fifo_csv_dumper_624,fifo_intf_624,cstatus_csv_dumper_624);
    fifo_csv_dumper_625 = new("./depth625.csv");
    cstatus_csv_dumper_625 = new("./chan_status625.csv");
    fifo_monitor_625 = new(fifo_csv_dumper_625,fifo_intf_625,cstatus_csv_dumper_625);
    fifo_csv_dumper_626 = new("./depth626.csv");
    cstatus_csv_dumper_626 = new("./chan_status626.csv");
    fifo_monitor_626 = new(fifo_csv_dumper_626,fifo_intf_626,cstatus_csv_dumper_626);
    fifo_csv_dumper_627 = new("./depth627.csv");
    cstatus_csv_dumper_627 = new("./chan_status627.csv");
    fifo_monitor_627 = new(fifo_csv_dumper_627,fifo_intf_627,cstatus_csv_dumper_627);
    fifo_csv_dumper_628 = new("./depth628.csv");
    cstatus_csv_dumper_628 = new("./chan_status628.csv");
    fifo_monitor_628 = new(fifo_csv_dumper_628,fifo_intf_628,cstatus_csv_dumper_628);
    fifo_csv_dumper_629 = new("./depth629.csv");
    cstatus_csv_dumper_629 = new("./chan_status629.csv");
    fifo_monitor_629 = new(fifo_csv_dumper_629,fifo_intf_629,cstatus_csv_dumper_629);
    fifo_csv_dumper_630 = new("./depth630.csv");
    cstatus_csv_dumper_630 = new("./chan_status630.csv");
    fifo_monitor_630 = new(fifo_csv_dumper_630,fifo_intf_630,cstatus_csv_dumper_630);
    fifo_csv_dumper_631 = new("./depth631.csv");
    cstatus_csv_dumper_631 = new("./chan_status631.csv");
    fifo_monitor_631 = new(fifo_csv_dumper_631,fifo_intf_631,cstatus_csv_dumper_631);
    fifo_csv_dumper_632 = new("./depth632.csv");
    cstatus_csv_dumper_632 = new("./chan_status632.csv");
    fifo_monitor_632 = new(fifo_csv_dumper_632,fifo_intf_632,cstatus_csv_dumper_632);
    fifo_csv_dumper_633 = new("./depth633.csv");
    cstatus_csv_dumper_633 = new("./chan_status633.csv");
    fifo_monitor_633 = new(fifo_csv_dumper_633,fifo_intf_633,cstatus_csv_dumper_633);
    fifo_csv_dumper_634 = new("./depth634.csv");
    cstatus_csv_dumper_634 = new("./chan_status634.csv");
    fifo_monitor_634 = new(fifo_csv_dumper_634,fifo_intf_634,cstatus_csv_dumper_634);
    fifo_csv_dumper_635 = new("./depth635.csv");
    cstatus_csv_dumper_635 = new("./chan_status635.csv");
    fifo_monitor_635 = new(fifo_csv_dumper_635,fifo_intf_635,cstatus_csv_dumper_635);
    fifo_csv_dumper_636 = new("./depth636.csv");
    cstatus_csv_dumper_636 = new("./chan_status636.csv");
    fifo_monitor_636 = new(fifo_csv_dumper_636,fifo_intf_636,cstatus_csv_dumper_636);
    fifo_csv_dumper_637 = new("./depth637.csv");
    cstatus_csv_dumper_637 = new("./chan_status637.csv");
    fifo_monitor_637 = new(fifo_csv_dumper_637,fifo_intf_637,cstatus_csv_dumper_637);
    fifo_csv_dumper_638 = new("./depth638.csv");
    cstatus_csv_dumper_638 = new("./chan_status638.csv");
    fifo_monitor_638 = new(fifo_csv_dumper_638,fifo_intf_638,cstatus_csv_dumper_638);
    fifo_csv_dumper_639 = new("./depth639.csv");
    cstatus_csv_dumper_639 = new("./chan_status639.csv");
    fifo_monitor_639 = new(fifo_csv_dumper_639,fifo_intf_639,cstatus_csv_dumper_639);
    fifo_csv_dumper_640 = new("./depth640.csv");
    cstatus_csv_dumper_640 = new("./chan_status640.csv");
    fifo_monitor_640 = new(fifo_csv_dumper_640,fifo_intf_640,cstatus_csv_dumper_640);
    fifo_csv_dumper_641 = new("./depth641.csv");
    cstatus_csv_dumper_641 = new("./chan_status641.csv");
    fifo_monitor_641 = new(fifo_csv_dumper_641,fifo_intf_641,cstatus_csv_dumper_641);
    fifo_csv_dumper_642 = new("./depth642.csv");
    cstatus_csv_dumper_642 = new("./chan_status642.csv");
    fifo_monitor_642 = new(fifo_csv_dumper_642,fifo_intf_642,cstatus_csv_dumper_642);
    fifo_csv_dumper_643 = new("./depth643.csv");
    cstatus_csv_dumper_643 = new("./chan_status643.csv");
    fifo_monitor_643 = new(fifo_csv_dumper_643,fifo_intf_643,cstatus_csv_dumper_643);
    fifo_csv_dumper_644 = new("./depth644.csv");
    cstatus_csv_dumper_644 = new("./chan_status644.csv");
    fifo_monitor_644 = new(fifo_csv_dumper_644,fifo_intf_644,cstatus_csv_dumper_644);
    fifo_csv_dumper_645 = new("./depth645.csv");
    cstatus_csv_dumper_645 = new("./chan_status645.csv");
    fifo_monitor_645 = new(fifo_csv_dumper_645,fifo_intf_645,cstatus_csv_dumper_645);
    fifo_csv_dumper_646 = new("./depth646.csv");
    cstatus_csv_dumper_646 = new("./chan_status646.csv");
    fifo_monitor_646 = new(fifo_csv_dumper_646,fifo_intf_646,cstatus_csv_dumper_646);
    fifo_csv_dumper_647 = new("./depth647.csv");
    cstatus_csv_dumper_647 = new("./chan_status647.csv");
    fifo_monitor_647 = new(fifo_csv_dumper_647,fifo_intf_647,cstatus_csv_dumper_647);
    fifo_csv_dumper_648 = new("./depth648.csv");
    cstatus_csv_dumper_648 = new("./chan_status648.csv");
    fifo_monitor_648 = new(fifo_csv_dumper_648,fifo_intf_648,cstatus_csv_dumper_648);
    fifo_csv_dumper_649 = new("./depth649.csv");
    cstatus_csv_dumper_649 = new("./chan_status649.csv");
    fifo_monitor_649 = new(fifo_csv_dumper_649,fifo_intf_649,cstatus_csv_dumper_649);
    fifo_csv_dumper_650 = new("./depth650.csv");
    cstatus_csv_dumper_650 = new("./chan_status650.csv");
    fifo_monitor_650 = new(fifo_csv_dumper_650,fifo_intf_650,cstatus_csv_dumper_650);
    fifo_csv_dumper_651 = new("./depth651.csv");
    cstatus_csv_dumper_651 = new("./chan_status651.csv");
    fifo_monitor_651 = new(fifo_csv_dumper_651,fifo_intf_651,cstatus_csv_dumper_651);
    fifo_csv_dumper_652 = new("./depth652.csv");
    cstatus_csv_dumper_652 = new("./chan_status652.csv");
    fifo_monitor_652 = new(fifo_csv_dumper_652,fifo_intf_652,cstatus_csv_dumper_652);
    fifo_csv_dumper_653 = new("./depth653.csv");
    cstatus_csv_dumper_653 = new("./chan_status653.csv");
    fifo_monitor_653 = new(fifo_csv_dumper_653,fifo_intf_653,cstatus_csv_dumper_653);
    fifo_csv_dumper_654 = new("./depth654.csv");
    cstatus_csv_dumper_654 = new("./chan_status654.csv");
    fifo_monitor_654 = new(fifo_csv_dumper_654,fifo_intf_654,cstatus_csv_dumper_654);
    fifo_csv_dumper_655 = new("./depth655.csv");
    cstatus_csv_dumper_655 = new("./chan_status655.csv");
    fifo_monitor_655 = new(fifo_csv_dumper_655,fifo_intf_655,cstatus_csv_dumper_655);
    fifo_csv_dumper_656 = new("./depth656.csv");
    cstatus_csv_dumper_656 = new("./chan_status656.csv");
    fifo_monitor_656 = new(fifo_csv_dumper_656,fifo_intf_656,cstatus_csv_dumper_656);
    fifo_csv_dumper_657 = new("./depth657.csv");
    cstatus_csv_dumper_657 = new("./chan_status657.csv");
    fifo_monitor_657 = new(fifo_csv_dumper_657,fifo_intf_657,cstatus_csv_dumper_657);
    fifo_csv_dumper_658 = new("./depth658.csv");
    cstatus_csv_dumper_658 = new("./chan_status658.csv");
    fifo_monitor_658 = new(fifo_csv_dumper_658,fifo_intf_658,cstatus_csv_dumper_658);
    fifo_csv_dumper_659 = new("./depth659.csv");
    cstatus_csv_dumper_659 = new("./chan_status659.csv");
    fifo_monitor_659 = new(fifo_csv_dumper_659,fifo_intf_659,cstatus_csv_dumper_659);
    fifo_csv_dumper_660 = new("./depth660.csv");
    cstatus_csv_dumper_660 = new("./chan_status660.csv");
    fifo_monitor_660 = new(fifo_csv_dumper_660,fifo_intf_660,cstatus_csv_dumper_660);
    fifo_csv_dumper_661 = new("./depth661.csv");
    cstatus_csv_dumper_661 = new("./chan_status661.csv");
    fifo_monitor_661 = new(fifo_csv_dumper_661,fifo_intf_661,cstatus_csv_dumper_661);
    fifo_csv_dumper_662 = new("./depth662.csv");
    cstatus_csv_dumper_662 = new("./chan_status662.csv");
    fifo_monitor_662 = new(fifo_csv_dumper_662,fifo_intf_662,cstatus_csv_dumper_662);
    fifo_csv_dumper_663 = new("./depth663.csv");
    cstatus_csv_dumper_663 = new("./chan_status663.csv");
    fifo_monitor_663 = new(fifo_csv_dumper_663,fifo_intf_663,cstatus_csv_dumper_663);
    fifo_csv_dumper_664 = new("./depth664.csv");
    cstatus_csv_dumper_664 = new("./chan_status664.csv");
    fifo_monitor_664 = new(fifo_csv_dumper_664,fifo_intf_664,cstatus_csv_dumper_664);
    fifo_csv_dumper_665 = new("./depth665.csv");
    cstatus_csv_dumper_665 = new("./chan_status665.csv");
    fifo_monitor_665 = new(fifo_csv_dumper_665,fifo_intf_665,cstatus_csv_dumper_665);
    fifo_csv_dumper_666 = new("./depth666.csv");
    cstatus_csv_dumper_666 = new("./chan_status666.csv");
    fifo_monitor_666 = new(fifo_csv_dumper_666,fifo_intf_666,cstatus_csv_dumper_666);
    fifo_csv_dumper_667 = new("./depth667.csv");
    cstatus_csv_dumper_667 = new("./chan_status667.csv");
    fifo_monitor_667 = new(fifo_csv_dumper_667,fifo_intf_667,cstatus_csv_dumper_667);
    fifo_csv_dumper_668 = new("./depth668.csv");
    cstatus_csv_dumper_668 = new("./chan_status668.csv");
    fifo_monitor_668 = new(fifo_csv_dumper_668,fifo_intf_668,cstatus_csv_dumper_668);
    fifo_csv_dumper_669 = new("./depth669.csv");
    cstatus_csv_dumper_669 = new("./chan_status669.csv");
    fifo_monitor_669 = new(fifo_csv_dumper_669,fifo_intf_669,cstatus_csv_dumper_669);
    fifo_csv_dumper_670 = new("./depth670.csv");
    cstatus_csv_dumper_670 = new("./chan_status670.csv");
    fifo_monitor_670 = new(fifo_csv_dumper_670,fifo_intf_670,cstatus_csv_dumper_670);
    fifo_csv_dumper_671 = new("./depth671.csv");
    cstatus_csv_dumper_671 = new("./chan_status671.csv");
    fifo_monitor_671 = new(fifo_csv_dumper_671,fifo_intf_671,cstatus_csv_dumper_671);
    fifo_csv_dumper_672 = new("./depth672.csv");
    cstatus_csv_dumper_672 = new("./chan_status672.csv");
    fifo_monitor_672 = new(fifo_csv_dumper_672,fifo_intf_672,cstatus_csv_dumper_672);
    fifo_csv_dumper_673 = new("./depth673.csv");
    cstatus_csv_dumper_673 = new("./chan_status673.csv");
    fifo_monitor_673 = new(fifo_csv_dumper_673,fifo_intf_673,cstatus_csv_dumper_673);
    fifo_csv_dumper_674 = new("./depth674.csv");
    cstatus_csv_dumper_674 = new("./chan_status674.csv");
    fifo_monitor_674 = new(fifo_csv_dumper_674,fifo_intf_674,cstatus_csv_dumper_674);
    fifo_csv_dumper_675 = new("./depth675.csv");
    cstatus_csv_dumper_675 = new("./chan_status675.csv");
    fifo_monitor_675 = new(fifo_csv_dumper_675,fifo_intf_675,cstatus_csv_dumper_675);
    fifo_csv_dumper_676 = new("./depth676.csv");
    cstatus_csv_dumper_676 = new("./chan_status676.csv");
    fifo_monitor_676 = new(fifo_csv_dumper_676,fifo_intf_676,cstatus_csv_dumper_676);
    fifo_csv_dumper_677 = new("./depth677.csv");
    cstatus_csv_dumper_677 = new("./chan_status677.csv");
    fifo_monitor_677 = new(fifo_csv_dumper_677,fifo_intf_677,cstatus_csv_dumper_677);
    fifo_csv_dumper_678 = new("./depth678.csv");
    cstatus_csv_dumper_678 = new("./chan_status678.csv");
    fifo_monitor_678 = new(fifo_csv_dumper_678,fifo_intf_678,cstatus_csv_dumper_678);
    fifo_csv_dumper_679 = new("./depth679.csv");
    cstatus_csv_dumper_679 = new("./chan_status679.csv");
    fifo_monitor_679 = new(fifo_csv_dumper_679,fifo_intf_679,cstatus_csv_dumper_679);
    fifo_csv_dumper_680 = new("./depth680.csv");
    cstatus_csv_dumper_680 = new("./chan_status680.csv");
    fifo_monitor_680 = new(fifo_csv_dumper_680,fifo_intf_680,cstatus_csv_dumper_680);
    fifo_csv_dumper_681 = new("./depth681.csv");
    cstatus_csv_dumper_681 = new("./chan_status681.csv");
    fifo_monitor_681 = new(fifo_csv_dumper_681,fifo_intf_681,cstatus_csv_dumper_681);
    fifo_csv_dumper_682 = new("./depth682.csv");
    cstatus_csv_dumper_682 = new("./chan_status682.csv");
    fifo_monitor_682 = new(fifo_csv_dumper_682,fifo_intf_682,cstatus_csv_dumper_682);
    fifo_csv_dumper_683 = new("./depth683.csv");
    cstatus_csv_dumper_683 = new("./chan_status683.csv");
    fifo_monitor_683 = new(fifo_csv_dumper_683,fifo_intf_683,cstatus_csv_dumper_683);
    fifo_csv_dumper_684 = new("./depth684.csv");
    cstatus_csv_dumper_684 = new("./chan_status684.csv");
    fifo_monitor_684 = new(fifo_csv_dumper_684,fifo_intf_684,cstatus_csv_dumper_684);
    fifo_csv_dumper_685 = new("./depth685.csv");
    cstatus_csv_dumper_685 = new("./chan_status685.csv");
    fifo_monitor_685 = new(fifo_csv_dumper_685,fifo_intf_685,cstatus_csv_dumper_685);
    fifo_csv_dumper_686 = new("./depth686.csv");
    cstatus_csv_dumper_686 = new("./chan_status686.csv");
    fifo_monitor_686 = new(fifo_csv_dumper_686,fifo_intf_686,cstatus_csv_dumper_686);
    fifo_csv_dumper_687 = new("./depth687.csv");
    cstatus_csv_dumper_687 = new("./chan_status687.csv");
    fifo_monitor_687 = new(fifo_csv_dumper_687,fifo_intf_687,cstatus_csv_dumper_687);
    fifo_csv_dumper_688 = new("./depth688.csv");
    cstatus_csv_dumper_688 = new("./chan_status688.csv");
    fifo_monitor_688 = new(fifo_csv_dumper_688,fifo_intf_688,cstatus_csv_dumper_688);
    fifo_csv_dumper_689 = new("./depth689.csv");
    cstatus_csv_dumper_689 = new("./chan_status689.csv");
    fifo_monitor_689 = new(fifo_csv_dumper_689,fifo_intf_689,cstatus_csv_dumper_689);
    fifo_csv_dumper_690 = new("./depth690.csv");
    cstatus_csv_dumper_690 = new("./chan_status690.csv");
    fifo_monitor_690 = new(fifo_csv_dumper_690,fifo_intf_690,cstatus_csv_dumper_690);
    fifo_csv_dumper_691 = new("./depth691.csv");
    cstatus_csv_dumper_691 = new("./chan_status691.csv");
    fifo_monitor_691 = new(fifo_csv_dumper_691,fifo_intf_691,cstatus_csv_dumper_691);
    fifo_csv_dumper_692 = new("./depth692.csv");
    cstatus_csv_dumper_692 = new("./chan_status692.csv");
    fifo_monitor_692 = new(fifo_csv_dumper_692,fifo_intf_692,cstatus_csv_dumper_692);
    fifo_csv_dumper_693 = new("./depth693.csv");
    cstatus_csv_dumper_693 = new("./chan_status693.csv");
    fifo_monitor_693 = new(fifo_csv_dumper_693,fifo_intf_693,cstatus_csv_dumper_693);
    fifo_csv_dumper_694 = new("./depth694.csv");
    cstatus_csv_dumper_694 = new("./chan_status694.csv");
    fifo_monitor_694 = new(fifo_csv_dumper_694,fifo_intf_694,cstatus_csv_dumper_694);
    fifo_csv_dumper_695 = new("./depth695.csv");
    cstatus_csv_dumper_695 = new("./chan_status695.csv");
    fifo_monitor_695 = new(fifo_csv_dumper_695,fifo_intf_695,cstatus_csv_dumper_695);
    fifo_csv_dumper_696 = new("./depth696.csv");
    cstatus_csv_dumper_696 = new("./chan_status696.csv");
    fifo_monitor_696 = new(fifo_csv_dumper_696,fifo_intf_696,cstatus_csv_dumper_696);
    fifo_csv_dumper_697 = new("./depth697.csv");
    cstatus_csv_dumper_697 = new("./chan_status697.csv");
    fifo_monitor_697 = new(fifo_csv_dumper_697,fifo_intf_697,cstatus_csv_dumper_697);
    fifo_csv_dumper_698 = new("./depth698.csv");
    cstatus_csv_dumper_698 = new("./chan_status698.csv");
    fifo_monitor_698 = new(fifo_csv_dumper_698,fifo_intf_698,cstatus_csv_dumper_698);
    fifo_csv_dumper_699 = new("./depth699.csv");
    cstatus_csv_dumper_699 = new("./chan_status699.csv");
    fifo_monitor_699 = new(fifo_csv_dumper_699,fifo_intf_699,cstatus_csv_dumper_699);
    fifo_csv_dumper_700 = new("./depth700.csv");
    cstatus_csv_dumper_700 = new("./chan_status700.csv");
    fifo_monitor_700 = new(fifo_csv_dumper_700,fifo_intf_700,cstatus_csv_dumper_700);
    fifo_csv_dumper_701 = new("./depth701.csv");
    cstatus_csv_dumper_701 = new("./chan_status701.csv");
    fifo_monitor_701 = new(fifo_csv_dumper_701,fifo_intf_701,cstatus_csv_dumper_701);
    fifo_csv_dumper_702 = new("./depth702.csv");
    cstatus_csv_dumper_702 = new("./chan_status702.csv");
    fifo_monitor_702 = new(fifo_csv_dumper_702,fifo_intf_702,cstatus_csv_dumper_702);
    fifo_csv_dumper_703 = new("./depth703.csv");
    cstatus_csv_dumper_703 = new("./chan_status703.csv");
    fifo_monitor_703 = new(fifo_csv_dumper_703,fifo_intf_703,cstatus_csv_dumper_703);
    fifo_csv_dumper_704 = new("./depth704.csv");
    cstatus_csv_dumper_704 = new("./chan_status704.csv");
    fifo_monitor_704 = new(fifo_csv_dumper_704,fifo_intf_704,cstatus_csv_dumper_704);
    fifo_csv_dumper_705 = new("./depth705.csv");
    cstatus_csv_dumper_705 = new("./chan_status705.csv");
    fifo_monitor_705 = new(fifo_csv_dumper_705,fifo_intf_705,cstatus_csv_dumper_705);
    fifo_csv_dumper_706 = new("./depth706.csv");
    cstatus_csv_dumper_706 = new("./chan_status706.csv");
    fifo_monitor_706 = new(fifo_csv_dumper_706,fifo_intf_706,cstatus_csv_dumper_706);
    fifo_csv_dumper_707 = new("./depth707.csv");
    cstatus_csv_dumper_707 = new("./chan_status707.csv");
    fifo_monitor_707 = new(fifo_csv_dumper_707,fifo_intf_707,cstatus_csv_dumper_707);
    fifo_csv_dumper_708 = new("./depth708.csv");
    cstatus_csv_dumper_708 = new("./chan_status708.csv");
    fifo_monitor_708 = new(fifo_csv_dumper_708,fifo_intf_708,cstatus_csv_dumper_708);
    fifo_csv_dumper_709 = new("./depth709.csv");
    cstatus_csv_dumper_709 = new("./chan_status709.csv");
    fifo_monitor_709 = new(fifo_csv_dumper_709,fifo_intf_709,cstatus_csv_dumper_709);
    fifo_csv_dumper_710 = new("./depth710.csv");
    cstatus_csv_dumper_710 = new("./chan_status710.csv");
    fifo_monitor_710 = new(fifo_csv_dumper_710,fifo_intf_710,cstatus_csv_dumper_710);
    fifo_csv_dumper_711 = new("./depth711.csv");
    cstatus_csv_dumper_711 = new("./chan_status711.csv");
    fifo_monitor_711 = new(fifo_csv_dumper_711,fifo_intf_711,cstatus_csv_dumper_711);
    fifo_csv_dumper_712 = new("./depth712.csv");
    cstatus_csv_dumper_712 = new("./chan_status712.csv");
    fifo_monitor_712 = new(fifo_csv_dumper_712,fifo_intf_712,cstatus_csv_dumper_712);
    fifo_csv_dumper_713 = new("./depth713.csv");
    cstatus_csv_dumper_713 = new("./chan_status713.csv");
    fifo_monitor_713 = new(fifo_csv_dumper_713,fifo_intf_713,cstatus_csv_dumper_713);
    fifo_csv_dumper_714 = new("./depth714.csv");
    cstatus_csv_dumper_714 = new("./chan_status714.csv");
    fifo_monitor_714 = new(fifo_csv_dumper_714,fifo_intf_714,cstatus_csv_dumper_714);
    fifo_csv_dumper_715 = new("./depth715.csv");
    cstatus_csv_dumper_715 = new("./chan_status715.csv");
    fifo_monitor_715 = new(fifo_csv_dumper_715,fifo_intf_715,cstatus_csv_dumper_715);
    fifo_csv_dumper_716 = new("./depth716.csv");
    cstatus_csv_dumper_716 = new("./chan_status716.csv");
    fifo_monitor_716 = new(fifo_csv_dumper_716,fifo_intf_716,cstatus_csv_dumper_716);
    fifo_csv_dumper_717 = new("./depth717.csv");
    cstatus_csv_dumper_717 = new("./chan_status717.csv");
    fifo_monitor_717 = new(fifo_csv_dumper_717,fifo_intf_717,cstatus_csv_dumper_717);
    fifo_csv_dumper_718 = new("./depth718.csv");
    cstatus_csv_dumper_718 = new("./chan_status718.csv");
    fifo_monitor_718 = new(fifo_csv_dumper_718,fifo_intf_718,cstatus_csv_dumper_718);
    fifo_csv_dumper_719 = new("./depth719.csv");
    cstatus_csv_dumper_719 = new("./chan_status719.csv");
    fifo_monitor_719 = new(fifo_csv_dumper_719,fifo_intf_719,cstatus_csv_dumper_719);
    fifo_csv_dumper_720 = new("./depth720.csv");
    cstatus_csv_dumper_720 = new("./chan_status720.csv");
    fifo_monitor_720 = new(fifo_csv_dumper_720,fifo_intf_720,cstatus_csv_dumper_720);
    fifo_csv_dumper_721 = new("./depth721.csv");
    cstatus_csv_dumper_721 = new("./chan_status721.csv");
    fifo_monitor_721 = new(fifo_csv_dumper_721,fifo_intf_721,cstatus_csv_dumper_721);
    fifo_csv_dumper_722 = new("./depth722.csv");
    cstatus_csv_dumper_722 = new("./chan_status722.csv");
    fifo_monitor_722 = new(fifo_csv_dumper_722,fifo_intf_722,cstatus_csv_dumper_722);
    fifo_csv_dumper_723 = new("./depth723.csv");
    cstatus_csv_dumper_723 = new("./chan_status723.csv");
    fifo_monitor_723 = new(fifo_csv_dumper_723,fifo_intf_723,cstatus_csv_dumper_723);
    fifo_csv_dumper_724 = new("./depth724.csv");
    cstatus_csv_dumper_724 = new("./chan_status724.csv");
    fifo_monitor_724 = new(fifo_csv_dumper_724,fifo_intf_724,cstatus_csv_dumper_724);
    fifo_csv_dumper_725 = new("./depth725.csv");
    cstatus_csv_dumper_725 = new("./chan_status725.csv");
    fifo_monitor_725 = new(fifo_csv_dumper_725,fifo_intf_725,cstatus_csv_dumper_725);
    fifo_csv_dumper_726 = new("./depth726.csv");
    cstatus_csv_dumper_726 = new("./chan_status726.csv");
    fifo_monitor_726 = new(fifo_csv_dumper_726,fifo_intf_726,cstatus_csv_dumper_726);
    fifo_csv_dumper_727 = new("./depth727.csv");
    cstatus_csv_dumper_727 = new("./chan_status727.csv");
    fifo_monitor_727 = new(fifo_csv_dumper_727,fifo_intf_727,cstatus_csv_dumper_727);
    fifo_csv_dumper_728 = new("./depth728.csv");
    cstatus_csv_dumper_728 = new("./chan_status728.csv");
    fifo_monitor_728 = new(fifo_csv_dumper_728,fifo_intf_728,cstatus_csv_dumper_728);
    fifo_csv_dumper_729 = new("./depth729.csv");
    cstatus_csv_dumper_729 = new("./chan_status729.csv");
    fifo_monitor_729 = new(fifo_csv_dumper_729,fifo_intf_729,cstatus_csv_dumper_729);
    fifo_csv_dumper_730 = new("./depth730.csv");
    cstatus_csv_dumper_730 = new("./chan_status730.csv");
    fifo_monitor_730 = new(fifo_csv_dumper_730,fifo_intf_730,cstatus_csv_dumper_730);
    fifo_csv_dumper_731 = new("./depth731.csv");
    cstatus_csv_dumper_731 = new("./chan_status731.csv");
    fifo_monitor_731 = new(fifo_csv_dumper_731,fifo_intf_731,cstatus_csv_dumper_731);
    fifo_csv_dumper_732 = new("./depth732.csv");
    cstatus_csv_dumper_732 = new("./chan_status732.csv");
    fifo_monitor_732 = new(fifo_csv_dumper_732,fifo_intf_732,cstatus_csv_dumper_732);
    fifo_csv_dumper_733 = new("./depth733.csv");
    cstatus_csv_dumper_733 = new("./chan_status733.csv");
    fifo_monitor_733 = new(fifo_csv_dumper_733,fifo_intf_733,cstatus_csv_dumper_733);
    fifo_csv_dumper_734 = new("./depth734.csv");
    cstatus_csv_dumper_734 = new("./chan_status734.csv");
    fifo_monitor_734 = new(fifo_csv_dumper_734,fifo_intf_734,cstatus_csv_dumper_734);
    fifo_csv_dumper_735 = new("./depth735.csv");
    cstatus_csv_dumper_735 = new("./chan_status735.csv");
    fifo_monitor_735 = new(fifo_csv_dumper_735,fifo_intf_735,cstatus_csv_dumper_735);
    fifo_csv_dumper_736 = new("./depth736.csv");
    cstatus_csv_dumper_736 = new("./chan_status736.csv");
    fifo_monitor_736 = new(fifo_csv_dumper_736,fifo_intf_736,cstatus_csv_dumper_736);
    fifo_csv_dumper_737 = new("./depth737.csv");
    cstatus_csv_dumper_737 = new("./chan_status737.csv");
    fifo_monitor_737 = new(fifo_csv_dumper_737,fifo_intf_737,cstatus_csv_dumper_737);
    fifo_csv_dumper_738 = new("./depth738.csv");
    cstatus_csv_dumper_738 = new("./chan_status738.csv");
    fifo_monitor_738 = new(fifo_csv_dumper_738,fifo_intf_738,cstatus_csv_dumper_738);
    fifo_csv_dumper_739 = new("./depth739.csv");
    cstatus_csv_dumper_739 = new("./chan_status739.csv");
    fifo_monitor_739 = new(fifo_csv_dumper_739,fifo_intf_739,cstatus_csv_dumper_739);
    fifo_csv_dumper_740 = new("./depth740.csv");
    cstatus_csv_dumper_740 = new("./chan_status740.csv");
    fifo_monitor_740 = new(fifo_csv_dumper_740,fifo_intf_740,cstatus_csv_dumper_740);
    fifo_csv_dumper_741 = new("./depth741.csv");
    cstatus_csv_dumper_741 = new("./chan_status741.csv");
    fifo_monitor_741 = new(fifo_csv_dumper_741,fifo_intf_741,cstatus_csv_dumper_741);
    fifo_csv_dumper_742 = new("./depth742.csv");
    cstatus_csv_dumper_742 = new("./chan_status742.csv");
    fifo_monitor_742 = new(fifo_csv_dumper_742,fifo_intf_742,cstatus_csv_dumper_742);
    fifo_csv_dumper_743 = new("./depth743.csv");
    cstatus_csv_dumper_743 = new("./chan_status743.csv");
    fifo_monitor_743 = new(fifo_csv_dumper_743,fifo_intf_743,cstatus_csv_dumper_743);
    fifo_csv_dumper_744 = new("./depth744.csv");
    cstatus_csv_dumper_744 = new("./chan_status744.csv");
    fifo_monitor_744 = new(fifo_csv_dumper_744,fifo_intf_744,cstatus_csv_dumper_744);
    fifo_csv_dumper_745 = new("./depth745.csv");
    cstatus_csv_dumper_745 = new("./chan_status745.csv");
    fifo_monitor_745 = new(fifo_csv_dumper_745,fifo_intf_745,cstatus_csv_dumper_745);
    fifo_csv_dumper_746 = new("./depth746.csv");
    cstatus_csv_dumper_746 = new("./chan_status746.csv");
    fifo_monitor_746 = new(fifo_csv_dumper_746,fifo_intf_746,cstatus_csv_dumper_746);
    fifo_csv_dumper_747 = new("./depth747.csv");
    cstatus_csv_dumper_747 = new("./chan_status747.csv");
    fifo_monitor_747 = new(fifo_csv_dumper_747,fifo_intf_747,cstatus_csv_dumper_747);
    fifo_csv_dumper_748 = new("./depth748.csv");
    cstatus_csv_dumper_748 = new("./chan_status748.csv");
    fifo_monitor_748 = new(fifo_csv_dumper_748,fifo_intf_748,cstatus_csv_dumper_748);
    fifo_csv_dumper_749 = new("./depth749.csv");
    cstatus_csv_dumper_749 = new("./chan_status749.csv");
    fifo_monitor_749 = new(fifo_csv_dumper_749,fifo_intf_749,cstatus_csv_dumper_749);
    fifo_csv_dumper_750 = new("./depth750.csv");
    cstatus_csv_dumper_750 = new("./chan_status750.csv");
    fifo_monitor_750 = new(fifo_csv_dumper_750,fifo_intf_750,cstatus_csv_dumper_750);
    fifo_csv_dumper_751 = new("./depth751.csv");
    cstatus_csv_dumper_751 = new("./chan_status751.csv");
    fifo_monitor_751 = new(fifo_csv_dumper_751,fifo_intf_751,cstatus_csv_dumper_751);
    fifo_csv_dumper_752 = new("./depth752.csv");
    cstatus_csv_dumper_752 = new("./chan_status752.csv");
    fifo_monitor_752 = new(fifo_csv_dumper_752,fifo_intf_752,cstatus_csv_dumper_752);
    fifo_csv_dumper_753 = new("./depth753.csv");
    cstatus_csv_dumper_753 = new("./chan_status753.csv");
    fifo_monitor_753 = new(fifo_csv_dumper_753,fifo_intf_753,cstatus_csv_dumper_753);
    fifo_csv_dumper_754 = new("./depth754.csv");
    cstatus_csv_dumper_754 = new("./chan_status754.csv");
    fifo_monitor_754 = new(fifo_csv_dumper_754,fifo_intf_754,cstatus_csv_dumper_754);
    fifo_csv_dumper_755 = new("./depth755.csv");
    cstatus_csv_dumper_755 = new("./chan_status755.csv");
    fifo_monitor_755 = new(fifo_csv_dumper_755,fifo_intf_755,cstatus_csv_dumper_755);
    fifo_csv_dumper_756 = new("./depth756.csv");
    cstatus_csv_dumper_756 = new("./chan_status756.csv");
    fifo_monitor_756 = new(fifo_csv_dumper_756,fifo_intf_756,cstatus_csv_dumper_756);
    fifo_csv_dumper_757 = new("./depth757.csv");
    cstatus_csv_dumper_757 = new("./chan_status757.csv");
    fifo_monitor_757 = new(fifo_csv_dumper_757,fifo_intf_757,cstatus_csv_dumper_757);
    fifo_csv_dumper_758 = new("./depth758.csv");
    cstatus_csv_dumper_758 = new("./chan_status758.csv");
    fifo_monitor_758 = new(fifo_csv_dumper_758,fifo_intf_758,cstatus_csv_dumper_758);
    fifo_csv_dumper_759 = new("./depth759.csv");
    cstatus_csv_dumper_759 = new("./chan_status759.csv");
    fifo_monitor_759 = new(fifo_csv_dumper_759,fifo_intf_759,cstatus_csv_dumper_759);
    fifo_csv_dumper_760 = new("./depth760.csv");
    cstatus_csv_dumper_760 = new("./chan_status760.csv");
    fifo_monitor_760 = new(fifo_csv_dumper_760,fifo_intf_760,cstatus_csv_dumper_760);
    fifo_csv_dumper_761 = new("./depth761.csv");
    cstatus_csv_dumper_761 = new("./chan_status761.csv");
    fifo_monitor_761 = new(fifo_csv_dumper_761,fifo_intf_761,cstatus_csv_dumper_761);
    fifo_csv_dumper_762 = new("./depth762.csv");
    cstatus_csv_dumper_762 = new("./chan_status762.csv");
    fifo_monitor_762 = new(fifo_csv_dumper_762,fifo_intf_762,cstatus_csv_dumper_762);
    fifo_csv_dumper_763 = new("./depth763.csv");
    cstatus_csv_dumper_763 = new("./chan_status763.csv");
    fifo_monitor_763 = new(fifo_csv_dumper_763,fifo_intf_763,cstatus_csv_dumper_763);
    fifo_csv_dumper_764 = new("./depth764.csv");
    cstatus_csv_dumper_764 = new("./chan_status764.csv");
    fifo_monitor_764 = new(fifo_csv_dumper_764,fifo_intf_764,cstatus_csv_dumper_764);
    fifo_csv_dumper_765 = new("./depth765.csv");
    cstatus_csv_dumper_765 = new("./chan_status765.csv");
    fifo_monitor_765 = new(fifo_csv_dumper_765,fifo_intf_765,cstatus_csv_dumper_765);
    fifo_csv_dumper_766 = new("./depth766.csv");
    cstatus_csv_dumper_766 = new("./chan_status766.csv");
    fifo_monitor_766 = new(fifo_csv_dumper_766,fifo_intf_766,cstatus_csv_dumper_766);
    fifo_csv_dumper_767 = new("./depth767.csv");
    cstatus_csv_dumper_767 = new("./chan_status767.csv");
    fifo_monitor_767 = new(fifo_csv_dumper_767,fifo_intf_767,cstatus_csv_dumper_767);
    fifo_csv_dumper_768 = new("./depth768.csv");
    cstatus_csv_dumper_768 = new("./chan_status768.csv");
    fifo_monitor_768 = new(fifo_csv_dumper_768,fifo_intf_768,cstatus_csv_dumper_768);
    fifo_csv_dumper_769 = new("./depth769.csv");
    cstatus_csv_dumper_769 = new("./chan_status769.csv");
    fifo_monitor_769 = new(fifo_csv_dumper_769,fifo_intf_769,cstatus_csv_dumper_769);
    fifo_csv_dumper_770 = new("./depth770.csv");
    cstatus_csv_dumper_770 = new("./chan_status770.csv");
    fifo_monitor_770 = new(fifo_csv_dumper_770,fifo_intf_770,cstatus_csv_dumper_770);
    fifo_csv_dumper_771 = new("./depth771.csv");
    cstatus_csv_dumper_771 = new("./chan_status771.csv");
    fifo_monitor_771 = new(fifo_csv_dumper_771,fifo_intf_771,cstatus_csv_dumper_771);
    fifo_csv_dumper_772 = new("./depth772.csv");
    cstatus_csv_dumper_772 = new("./chan_status772.csv");
    fifo_monitor_772 = new(fifo_csv_dumper_772,fifo_intf_772,cstatus_csv_dumper_772);
    fifo_csv_dumper_773 = new("./depth773.csv");
    cstatus_csv_dumper_773 = new("./chan_status773.csv");
    fifo_monitor_773 = new(fifo_csv_dumper_773,fifo_intf_773,cstatus_csv_dumper_773);
    fifo_csv_dumper_774 = new("./depth774.csv");
    cstatus_csv_dumper_774 = new("./chan_status774.csv");
    fifo_monitor_774 = new(fifo_csv_dumper_774,fifo_intf_774,cstatus_csv_dumper_774);
    fifo_csv_dumper_775 = new("./depth775.csv");
    cstatus_csv_dumper_775 = new("./chan_status775.csv");
    fifo_monitor_775 = new(fifo_csv_dumper_775,fifo_intf_775,cstatus_csv_dumper_775);
    fifo_csv_dumper_776 = new("./depth776.csv");
    cstatus_csv_dumper_776 = new("./chan_status776.csv");
    fifo_monitor_776 = new(fifo_csv_dumper_776,fifo_intf_776,cstatus_csv_dumper_776);
    fifo_csv_dumper_777 = new("./depth777.csv");
    cstatus_csv_dumper_777 = new("./chan_status777.csv");
    fifo_monitor_777 = new(fifo_csv_dumper_777,fifo_intf_777,cstatus_csv_dumper_777);
    fifo_csv_dumper_778 = new("./depth778.csv");
    cstatus_csv_dumper_778 = new("./chan_status778.csv");
    fifo_monitor_778 = new(fifo_csv_dumper_778,fifo_intf_778,cstatus_csv_dumper_778);
    fifo_csv_dumper_779 = new("./depth779.csv");
    cstatus_csv_dumper_779 = new("./chan_status779.csv");
    fifo_monitor_779 = new(fifo_csv_dumper_779,fifo_intf_779,cstatus_csv_dumper_779);
    fifo_csv_dumper_780 = new("./depth780.csv");
    cstatus_csv_dumper_780 = new("./chan_status780.csv");
    fifo_monitor_780 = new(fifo_csv_dumper_780,fifo_intf_780,cstatus_csv_dumper_780);
    fifo_csv_dumper_781 = new("./depth781.csv");
    cstatus_csv_dumper_781 = new("./chan_status781.csv");
    fifo_monitor_781 = new(fifo_csv_dumper_781,fifo_intf_781,cstatus_csv_dumper_781);
    fifo_csv_dumper_782 = new("./depth782.csv");
    cstatus_csv_dumper_782 = new("./chan_status782.csv");
    fifo_monitor_782 = new(fifo_csv_dumper_782,fifo_intf_782,cstatus_csv_dumper_782);
    fifo_csv_dumper_783 = new("./depth783.csv");
    cstatus_csv_dumper_783 = new("./chan_status783.csv");
    fifo_monitor_783 = new(fifo_csv_dumper_783,fifo_intf_783,cstatus_csv_dumper_783);
    fifo_csv_dumper_784 = new("./depth784.csv");
    cstatus_csv_dumper_784 = new("./chan_status784.csv");
    fifo_monitor_784 = new(fifo_csv_dumper_784,fifo_intf_784,cstatus_csv_dumper_784);
    fifo_csv_dumper_785 = new("./depth785.csv");
    cstatus_csv_dumper_785 = new("./chan_status785.csv");
    fifo_monitor_785 = new(fifo_csv_dumper_785,fifo_intf_785,cstatus_csv_dumper_785);
    fifo_csv_dumper_786 = new("./depth786.csv");
    cstatus_csv_dumper_786 = new("./chan_status786.csv");
    fifo_monitor_786 = new(fifo_csv_dumper_786,fifo_intf_786,cstatus_csv_dumper_786);
    fifo_csv_dumper_787 = new("./depth787.csv");
    cstatus_csv_dumper_787 = new("./chan_status787.csv");
    fifo_monitor_787 = new(fifo_csv_dumper_787,fifo_intf_787,cstatus_csv_dumper_787);
    fifo_csv_dumper_788 = new("./depth788.csv");
    cstatus_csv_dumper_788 = new("./chan_status788.csv");
    fifo_monitor_788 = new(fifo_csv_dumper_788,fifo_intf_788,cstatus_csv_dumper_788);
    fifo_csv_dumper_789 = new("./depth789.csv");
    cstatus_csv_dumper_789 = new("./chan_status789.csv");
    fifo_monitor_789 = new(fifo_csv_dumper_789,fifo_intf_789,cstatus_csv_dumper_789);
    fifo_csv_dumper_790 = new("./depth790.csv");
    cstatus_csv_dumper_790 = new("./chan_status790.csv");
    fifo_monitor_790 = new(fifo_csv_dumper_790,fifo_intf_790,cstatus_csv_dumper_790);
    fifo_csv_dumper_791 = new("./depth791.csv");
    cstatus_csv_dumper_791 = new("./chan_status791.csv");
    fifo_monitor_791 = new(fifo_csv_dumper_791,fifo_intf_791,cstatus_csv_dumper_791);
    fifo_csv_dumper_792 = new("./depth792.csv");
    cstatus_csv_dumper_792 = new("./chan_status792.csv");
    fifo_monitor_792 = new(fifo_csv_dumper_792,fifo_intf_792,cstatus_csv_dumper_792);
    fifo_csv_dumper_793 = new("./depth793.csv");
    cstatus_csv_dumper_793 = new("./chan_status793.csv");
    fifo_monitor_793 = new(fifo_csv_dumper_793,fifo_intf_793,cstatus_csv_dumper_793);
    fifo_csv_dumper_794 = new("./depth794.csv");
    cstatus_csv_dumper_794 = new("./chan_status794.csv");
    fifo_monitor_794 = new(fifo_csv_dumper_794,fifo_intf_794,cstatus_csv_dumper_794);
    fifo_csv_dumper_795 = new("./depth795.csv");
    cstatus_csv_dumper_795 = new("./chan_status795.csv");
    fifo_monitor_795 = new(fifo_csv_dumper_795,fifo_intf_795,cstatus_csv_dumper_795);
    fifo_csv_dumper_796 = new("./depth796.csv");
    cstatus_csv_dumper_796 = new("./chan_status796.csv");
    fifo_monitor_796 = new(fifo_csv_dumper_796,fifo_intf_796,cstatus_csv_dumper_796);
    fifo_csv_dumper_797 = new("./depth797.csv");
    cstatus_csv_dumper_797 = new("./chan_status797.csv");
    fifo_monitor_797 = new(fifo_csv_dumper_797,fifo_intf_797,cstatus_csv_dumper_797);
    fifo_csv_dumper_798 = new("./depth798.csv");
    cstatus_csv_dumper_798 = new("./chan_status798.csv");
    fifo_monitor_798 = new(fifo_csv_dumper_798,fifo_intf_798,cstatus_csv_dumper_798);
    fifo_csv_dumper_799 = new("./depth799.csv");
    cstatus_csv_dumper_799 = new("./chan_status799.csv");
    fifo_monitor_799 = new(fifo_csv_dumper_799,fifo_intf_799,cstatus_csv_dumper_799);
    fifo_csv_dumper_800 = new("./depth800.csv");
    cstatus_csv_dumper_800 = new("./chan_status800.csv");
    fifo_monitor_800 = new(fifo_csv_dumper_800,fifo_intf_800,cstatus_csv_dumper_800);
    fifo_csv_dumper_801 = new("./depth801.csv");
    cstatus_csv_dumper_801 = new("./chan_status801.csv");
    fifo_monitor_801 = new(fifo_csv_dumper_801,fifo_intf_801,cstatus_csv_dumper_801);
    fifo_csv_dumper_802 = new("./depth802.csv");
    cstatus_csv_dumper_802 = new("./chan_status802.csv");
    fifo_monitor_802 = new(fifo_csv_dumper_802,fifo_intf_802,cstatus_csv_dumper_802);
    fifo_csv_dumper_803 = new("./depth803.csv");
    cstatus_csv_dumper_803 = new("./chan_status803.csv");
    fifo_monitor_803 = new(fifo_csv_dumper_803,fifo_intf_803,cstatus_csv_dumper_803);
    fifo_csv_dumper_804 = new("./depth804.csv");
    cstatus_csv_dumper_804 = new("./chan_status804.csv");
    fifo_monitor_804 = new(fifo_csv_dumper_804,fifo_intf_804,cstatus_csv_dumper_804);
    fifo_csv_dumper_805 = new("./depth805.csv");
    cstatus_csv_dumper_805 = new("./chan_status805.csv");
    fifo_monitor_805 = new(fifo_csv_dumper_805,fifo_intf_805,cstatus_csv_dumper_805);
    fifo_csv_dumper_806 = new("./depth806.csv");
    cstatus_csv_dumper_806 = new("./chan_status806.csv");
    fifo_monitor_806 = new(fifo_csv_dumper_806,fifo_intf_806,cstatus_csv_dumper_806);
    fifo_csv_dumper_807 = new("./depth807.csv");
    cstatus_csv_dumper_807 = new("./chan_status807.csv");
    fifo_monitor_807 = new(fifo_csv_dumper_807,fifo_intf_807,cstatus_csv_dumper_807);
    fifo_csv_dumper_808 = new("./depth808.csv");
    cstatus_csv_dumper_808 = new("./chan_status808.csv");
    fifo_monitor_808 = new(fifo_csv_dumper_808,fifo_intf_808,cstatus_csv_dumper_808);
    fifo_csv_dumper_809 = new("./depth809.csv");
    cstatus_csv_dumper_809 = new("./chan_status809.csv");
    fifo_monitor_809 = new(fifo_csv_dumper_809,fifo_intf_809,cstatus_csv_dumper_809);
    fifo_csv_dumper_810 = new("./depth810.csv");
    cstatus_csv_dumper_810 = new("./chan_status810.csv");
    fifo_monitor_810 = new(fifo_csv_dumper_810,fifo_intf_810,cstatus_csv_dumper_810);
    fifo_csv_dumper_811 = new("./depth811.csv");
    cstatus_csv_dumper_811 = new("./chan_status811.csv");
    fifo_monitor_811 = new(fifo_csv_dumper_811,fifo_intf_811,cstatus_csv_dumper_811);
    fifo_csv_dumper_812 = new("./depth812.csv");
    cstatus_csv_dumper_812 = new("./chan_status812.csv");
    fifo_monitor_812 = new(fifo_csv_dumper_812,fifo_intf_812,cstatus_csv_dumper_812);
    fifo_csv_dumper_813 = new("./depth813.csv");
    cstatus_csv_dumper_813 = new("./chan_status813.csv");
    fifo_monitor_813 = new(fifo_csv_dumper_813,fifo_intf_813,cstatus_csv_dumper_813);
    fifo_csv_dumper_814 = new("./depth814.csv");
    cstatus_csv_dumper_814 = new("./chan_status814.csv");
    fifo_monitor_814 = new(fifo_csv_dumper_814,fifo_intf_814,cstatus_csv_dumper_814);
    fifo_csv_dumper_815 = new("./depth815.csv");
    cstatus_csv_dumper_815 = new("./chan_status815.csv");
    fifo_monitor_815 = new(fifo_csv_dumper_815,fifo_intf_815,cstatus_csv_dumper_815);
    fifo_csv_dumper_816 = new("./depth816.csv");
    cstatus_csv_dumper_816 = new("./chan_status816.csv");
    fifo_monitor_816 = new(fifo_csv_dumper_816,fifo_intf_816,cstatus_csv_dumper_816);
    fifo_csv_dumper_817 = new("./depth817.csv");
    cstatus_csv_dumper_817 = new("./chan_status817.csv");
    fifo_monitor_817 = new(fifo_csv_dumper_817,fifo_intf_817,cstatus_csv_dumper_817);
    fifo_csv_dumper_818 = new("./depth818.csv");
    cstatus_csv_dumper_818 = new("./chan_status818.csv");
    fifo_monitor_818 = new(fifo_csv_dumper_818,fifo_intf_818,cstatus_csv_dumper_818);
    fifo_csv_dumper_819 = new("./depth819.csv");
    cstatus_csv_dumper_819 = new("./chan_status819.csv");
    fifo_monitor_819 = new(fifo_csv_dumper_819,fifo_intf_819,cstatus_csv_dumper_819);
    fifo_csv_dumper_820 = new("./depth820.csv");
    cstatus_csv_dumper_820 = new("./chan_status820.csv");
    fifo_monitor_820 = new(fifo_csv_dumper_820,fifo_intf_820,cstatus_csv_dumper_820);
    fifo_csv_dumper_821 = new("./depth821.csv");
    cstatus_csv_dumper_821 = new("./chan_status821.csv");
    fifo_monitor_821 = new(fifo_csv_dumper_821,fifo_intf_821,cstatus_csv_dumper_821);
    fifo_csv_dumper_822 = new("./depth822.csv");
    cstatus_csv_dumper_822 = new("./chan_status822.csv");
    fifo_monitor_822 = new(fifo_csv_dumper_822,fifo_intf_822,cstatus_csv_dumper_822);
    fifo_csv_dumper_823 = new("./depth823.csv");
    cstatus_csv_dumper_823 = new("./chan_status823.csv");
    fifo_monitor_823 = new(fifo_csv_dumper_823,fifo_intf_823,cstatus_csv_dumper_823);
    fifo_csv_dumper_824 = new("./depth824.csv");
    cstatus_csv_dumper_824 = new("./chan_status824.csv");
    fifo_monitor_824 = new(fifo_csv_dumper_824,fifo_intf_824,cstatus_csv_dumper_824);
    fifo_csv_dumper_825 = new("./depth825.csv");
    cstatus_csv_dumper_825 = new("./chan_status825.csv");
    fifo_monitor_825 = new(fifo_csv_dumper_825,fifo_intf_825,cstatus_csv_dumper_825);
    fifo_csv_dumper_826 = new("./depth826.csv");
    cstatus_csv_dumper_826 = new("./chan_status826.csv");
    fifo_monitor_826 = new(fifo_csv_dumper_826,fifo_intf_826,cstatus_csv_dumper_826);
    fifo_csv_dumper_827 = new("./depth827.csv");
    cstatus_csv_dumper_827 = new("./chan_status827.csv");
    fifo_monitor_827 = new(fifo_csv_dumper_827,fifo_intf_827,cstatus_csv_dumper_827);
    fifo_csv_dumper_828 = new("./depth828.csv");
    cstatus_csv_dumper_828 = new("./chan_status828.csv");
    fifo_monitor_828 = new(fifo_csv_dumper_828,fifo_intf_828,cstatus_csv_dumper_828);
    fifo_csv_dumper_829 = new("./depth829.csv");
    cstatus_csv_dumper_829 = new("./chan_status829.csv");
    fifo_monitor_829 = new(fifo_csv_dumper_829,fifo_intf_829,cstatus_csv_dumper_829);
    fifo_csv_dumper_830 = new("./depth830.csv");
    cstatus_csv_dumper_830 = new("./chan_status830.csv");
    fifo_monitor_830 = new(fifo_csv_dumper_830,fifo_intf_830,cstatus_csv_dumper_830);
    fifo_csv_dumper_831 = new("./depth831.csv");
    cstatus_csv_dumper_831 = new("./chan_status831.csv");
    fifo_monitor_831 = new(fifo_csv_dumper_831,fifo_intf_831,cstatus_csv_dumper_831);
    fifo_csv_dumper_832 = new("./depth832.csv");
    cstatus_csv_dumper_832 = new("./chan_status832.csv");
    fifo_monitor_832 = new(fifo_csv_dumper_832,fifo_intf_832,cstatus_csv_dumper_832);
    fifo_csv_dumper_833 = new("./depth833.csv");
    cstatus_csv_dumper_833 = new("./chan_status833.csv");
    fifo_monitor_833 = new(fifo_csv_dumper_833,fifo_intf_833,cstatus_csv_dumper_833);
    fifo_csv_dumper_834 = new("./depth834.csv");
    cstatus_csv_dumper_834 = new("./chan_status834.csv");
    fifo_monitor_834 = new(fifo_csv_dumper_834,fifo_intf_834,cstatus_csv_dumper_834);
    fifo_csv_dumper_835 = new("./depth835.csv");
    cstatus_csv_dumper_835 = new("./chan_status835.csv");
    fifo_monitor_835 = new(fifo_csv_dumper_835,fifo_intf_835,cstatus_csv_dumper_835);
    fifo_csv_dumper_836 = new("./depth836.csv");
    cstatus_csv_dumper_836 = new("./chan_status836.csv");
    fifo_monitor_836 = new(fifo_csv_dumper_836,fifo_intf_836,cstatus_csv_dumper_836);
    fifo_csv_dumper_837 = new("./depth837.csv");
    cstatus_csv_dumper_837 = new("./chan_status837.csv");
    fifo_monitor_837 = new(fifo_csv_dumper_837,fifo_intf_837,cstatus_csv_dumper_837);
    fifo_csv_dumper_838 = new("./depth838.csv");
    cstatus_csv_dumper_838 = new("./chan_status838.csv");
    fifo_monitor_838 = new(fifo_csv_dumper_838,fifo_intf_838,cstatus_csv_dumper_838);
    fifo_csv_dumper_839 = new("./depth839.csv");
    cstatus_csv_dumper_839 = new("./chan_status839.csv");
    fifo_monitor_839 = new(fifo_csv_dumper_839,fifo_intf_839,cstatus_csv_dumper_839);
    fifo_csv_dumper_840 = new("./depth840.csv");
    cstatus_csv_dumper_840 = new("./chan_status840.csv");
    fifo_monitor_840 = new(fifo_csv_dumper_840,fifo_intf_840,cstatus_csv_dumper_840);
    fifo_csv_dumper_841 = new("./depth841.csv");
    cstatus_csv_dumper_841 = new("./chan_status841.csv");
    fifo_monitor_841 = new(fifo_csv_dumper_841,fifo_intf_841,cstatus_csv_dumper_841);
    fifo_csv_dumper_842 = new("./depth842.csv");
    cstatus_csv_dumper_842 = new("./chan_status842.csv");
    fifo_monitor_842 = new(fifo_csv_dumper_842,fifo_intf_842,cstatus_csv_dumper_842);
    fifo_csv_dumper_843 = new("./depth843.csv");
    cstatus_csv_dumper_843 = new("./chan_status843.csv");
    fifo_monitor_843 = new(fifo_csv_dumper_843,fifo_intf_843,cstatus_csv_dumper_843);
    fifo_csv_dumper_844 = new("./depth844.csv");
    cstatus_csv_dumper_844 = new("./chan_status844.csv");
    fifo_monitor_844 = new(fifo_csv_dumper_844,fifo_intf_844,cstatus_csv_dumper_844);
    fifo_csv_dumper_845 = new("./depth845.csv");
    cstatus_csv_dumper_845 = new("./chan_status845.csv");
    fifo_monitor_845 = new(fifo_csv_dumper_845,fifo_intf_845,cstatus_csv_dumper_845);
    fifo_csv_dumper_846 = new("./depth846.csv");
    cstatus_csv_dumper_846 = new("./chan_status846.csv");
    fifo_monitor_846 = new(fifo_csv_dumper_846,fifo_intf_846,cstatus_csv_dumper_846);
    fifo_csv_dumper_847 = new("./depth847.csv");
    cstatus_csv_dumper_847 = new("./chan_status847.csv");
    fifo_monitor_847 = new(fifo_csv_dumper_847,fifo_intf_847,cstatus_csv_dumper_847);
    fifo_csv_dumper_848 = new("./depth848.csv");
    cstatus_csv_dumper_848 = new("./chan_status848.csv");
    fifo_monitor_848 = new(fifo_csv_dumper_848,fifo_intf_848,cstatus_csv_dumper_848);
    fifo_csv_dumper_849 = new("./depth849.csv");
    cstatus_csv_dumper_849 = new("./chan_status849.csv");
    fifo_monitor_849 = new(fifo_csv_dumper_849,fifo_intf_849,cstatus_csv_dumper_849);
    fifo_csv_dumper_850 = new("./depth850.csv");
    cstatus_csv_dumper_850 = new("./chan_status850.csv");
    fifo_monitor_850 = new(fifo_csv_dumper_850,fifo_intf_850,cstatus_csv_dumper_850);
    fifo_csv_dumper_851 = new("./depth851.csv");
    cstatus_csv_dumper_851 = new("./chan_status851.csv");
    fifo_monitor_851 = new(fifo_csv_dumper_851,fifo_intf_851,cstatus_csv_dumper_851);
    fifo_csv_dumper_852 = new("./depth852.csv");
    cstatus_csv_dumper_852 = new("./chan_status852.csv");
    fifo_monitor_852 = new(fifo_csv_dumper_852,fifo_intf_852,cstatus_csv_dumper_852);
    fifo_csv_dumper_853 = new("./depth853.csv");
    cstatus_csv_dumper_853 = new("./chan_status853.csv");
    fifo_monitor_853 = new(fifo_csv_dumper_853,fifo_intf_853,cstatus_csv_dumper_853);
    fifo_csv_dumper_854 = new("./depth854.csv");
    cstatus_csv_dumper_854 = new("./chan_status854.csv");
    fifo_monitor_854 = new(fifo_csv_dumper_854,fifo_intf_854,cstatus_csv_dumper_854);
    fifo_csv_dumper_855 = new("./depth855.csv");
    cstatus_csv_dumper_855 = new("./chan_status855.csv");
    fifo_monitor_855 = new(fifo_csv_dumper_855,fifo_intf_855,cstatus_csv_dumper_855);
    fifo_csv_dumper_856 = new("./depth856.csv");
    cstatus_csv_dumper_856 = new("./chan_status856.csv");
    fifo_monitor_856 = new(fifo_csv_dumper_856,fifo_intf_856,cstatus_csv_dumper_856);
    fifo_csv_dumper_857 = new("./depth857.csv");
    cstatus_csv_dumper_857 = new("./chan_status857.csv");
    fifo_monitor_857 = new(fifo_csv_dumper_857,fifo_intf_857,cstatus_csv_dumper_857);
    fifo_csv_dumper_858 = new("./depth858.csv");
    cstatus_csv_dumper_858 = new("./chan_status858.csv");
    fifo_monitor_858 = new(fifo_csv_dumper_858,fifo_intf_858,cstatus_csv_dumper_858);
    fifo_csv_dumper_859 = new("./depth859.csv");
    cstatus_csv_dumper_859 = new("./chan_status859.csv");
    fifo_monitor_859 = new(fifo_csv_dumper_859,fifo_intf_859,cstatus_csv_dumper_859);
    fifo_csv_dumper_860 = new("./depth860.csv");
    cstatus_csv_dumper_860 = new("./chan_status860.csv");
    fifo_monitor_860 = new(fifo_csv_dumper_860,fifo_intf_860,cstatus_csv_dumper_860);
    fifo_csv_dumper_861 = new("./depth861.csv");
    cstatus_csv_dumper_861 = new("./chan_status861.csv");
    fifo_monitor_861 = new(fifo_csv_dumper_861,fifo_intf_861,cstatus_csv_dumper_861);
    fifo_csv_dumper_862 = new("./depth862.csv");
    cstatus_csv_dumper_862 = new("./chan_status862.csv");
    fifo_monitor_862 = new(fifo_csv_dumper_862,fifo_intf_862,cstatus_csv_dumper_862);
    fifo_csv_dumper_863 = new("./depth863.csv");
    cstatus_csv_dumper_863 = new("./chan_status863.csv");
    fifo_monitor_863 = new(fifo_csv_dumper_863,fifo_intf_863,cstatus_csv_dumper_863);
    fifo_csv_dumper_864 = new("./depth864.csv");
    cstatus_csv_dumper_864 = new("./chan_status864.csv");
    fifo_monitor_864 = new(fifo_csv_dumper_864,fifo_intf_864,cstatus_csv_dumper_864);
    fifo_csv_dumper_865 = new("./depth865.csv");
    cstatus_csv_dumper_865 = new("./chan_status865.csv");
    fifo_monitor_865 = new(fifo_csv_dumper_865,fifo_intf_865,cstatus_csv_dumper_865);
    fifo_csv_dumper_866 = new("./depth866.csv");
    cstatus_csv_dumper_866 = new("./chan_status866.csv");
    fifo_monitor_866 = new(fifo_csv_dumper_866,fifo_intf_866,cstatus_csv_dumper_866);
    fifo_csv_dumper_867 = new("./depth867.csv");
    cstatus_csv_dumper_867 = new("./chan_status867.csv");
    fifo_monitor_867 = new(fifo_csv_dumper_867,fifo_intf_867,cstatus_csv_dumper_867);
    fifo_csv_dumper_868 = new("./depth868.csv");
    cstatus_csv_dumper_868 = new("./chan_status868.csv");
    fifo_monitor_868 = new(fifo_csv_dumper_868,fifo_intf_868,cstatus_csv_dumper_868);
    fifo_csv_dumper_869 = new("./depth869.csv");
    cstatus_csv_dumper_869 = new("./chan_status869.csv");
    fifo_monitor_869 = new(fifo_csv_dumper_869,fifo_intf_869,cstatus_csv_dumper_869);
    fifo_csv_dumper_870 = new("./depth870.csv");
    cstatus_csv_dumper_870 = new("./chan_status870.csv");
    fifo_monitor_870 = new(fifo_csv_dumper_870,fifo_intf_870,cstatus_csv_dumper_870);
    fifo_csv_dumper_871 = new("./depth871.csv");
    cstatus_csv_dumper_871 = new("./chan_status871.csv");
    fifo_monitor_871 = new(fifo_csv_dumper_871,fifo_intf_871,cstatus_csv_dumper_871);
    fifo_csv_dumper_872 = new("./depth872.csv");
    cstatus_csv_dumper_872 = new("./chan_status872.csv");
    fifo_monitor_872 = new(fifo_csv_dumper_872,fifo_intf_872,cstatus_csv_dumper_872);
    fifo_csv_dumper_873 = new("./depth873.csv");
    cstatus_csv_dumper_873 = new("./chan_status873.csv");
    fifo_monitor_873 = new(fifo_csv_dumper_873,fifo_intf_873,cstatus_csv_dumper_873);
    fifo_csv_dumper_874 = new("./depth874.csv");
    cstatus_csv_dumper_874 = new("./chan_status874.csv");
    fifo_monitor_874 = new(fifo_csv_dumper_874,fifo_intf_874,cstatus_csv_dumper_874);
    fifo_csv_dumper_875 = new("./depth875.csv");
    cstatus_csv_dumper_875 = new("./chan_status875.csv");
    fifo_monitor_875 = new(fifo_csv_dumper_875,fifo_intf_875,cstatus_csv_dumper_875);
    fifo_csv_dumper_876 = new("./depth876.csv");
    cstatus_csv_dumper_876 = new("./chan_status876.csv");
    fifo_monitor_876 = new(fifo_csv_dumper_876,fifo_intf_876,cstatus_csv_dumper_876);
    fifo_csv_dumper_877 = new("./depth877.csv");
    cstatus_csv_dumper_877 = new("./chan_status877.csv");
    fifo_monitor_877 = new(fifo_csv_dumper_877,fifo_intf_877,cstatus_csv_dumper_877);
    fifo_csv_dumper_878 = new("./depth878.csv");
    cstatus_csv_dumper_878 = new("./chan_status878.csv");
    fifo_monitor_878 = new(fifo_csv_dumper_878,fifo_intf_878,cstatus_csv_dumper_878);
    fifo_csv_dumper_879 = new("./depth879.csv");
    cstatus_csv_dumper_879 = new("./chan_status879.csv");
    fifo_monitor_879 = new(fifo_csv_dumper_879,fifo_intf_879,cstatus_csv_dumper_879);
    fifo_csv_dumper_880 = new("./depth880.csv");
    cstatus_csv_dumper_880 = new("./chan_status880.csv");
    fifo_monitor_880 = new(fifo_csv_dumper_880,fifo_intf_880,cstatus_csv_dumper_880);
    fifo_csv_dumper_881 = new("./depth881.csv");
    cstatus_csv_dumper_881 = new("./chan_status881.csv");
    fifo_monitor_881 = new(fifo_csv_dumper_881,fifo_intf_881,cstatus_csv_dumper_881);
    fifo_csv_dumper_882 = new("./depth882.csv");
    cstatus_csv_dumper_882 = new("./chan_status882.csv");
    fifo_monitor_882 = new(fifo_csv_dumper_882,fifo_intf_882,cstatus_csv_dumper_882);
    fifo_csv_dumper_883 = new("./depth883.csv");
    cstatus_csv_dumper_883 = new("./chan_status883.csv");
    fifo_monitor_883 = new(fifo_csv_dumper_883,fifo_intf_883,cstatus_csv_dumper_883);
    fifo_csv_dumper_884 = new("./depth884.csv");
    cstatus_csv_dumper_884 = new("./chan_status884.csv");
    fifo_monitor_884 = new(fifo_csv_dumper_884,fifo_intf_884,cstatus_csv_dumper_884);
    fifo_csv_dumper_885 = new("./depth885.csv");
    cstatus_csv_dumper_885 = new("./chan_status885.csv");
    fifo_monitor_885 = new(fifo_csv_dumper_885,fifo_intf_885,cstatus_csv_dumper_885);
    fifo_csv_dumper_886 = new("./depth886.csv");
    cstatus_csv_dumper_886 = new("./chan_status886.csv");
    fifo_monitor_886 = new(fifo_csv_dumper_886,fifo_intf_886,cstatus_csv_dumper_886);
    fifo_csv_dumper_887 = new("./depth887.csv");
    cstatus_csv_dumper_887 = new("./chan_status887.csv");
    fifo_monitor_887 = new(fifo_csv_dumper_887,fifo_intf_887,cstatus_csv_dumper_887);
    fifo_csv_dumper_888 = new("./depth888.csv");
    cstatus_csv_dumper_888 = new("./chan_status888.csv");
    fifo_monitor_888 = new(fifo_csv_dumper_888,fifo_intf_888,cstatus_csv_dumper_888);
    fifo_csv_dumper_889 = new("./depth889.csv");
    cstatus_csv_dumper_889 = new("./chan_status889.csv");
    fifo_monitor_889 = new(fifo_csv_dumper_889,fifo_intf_889,cstatus_csv_dumper_889);
    fifo_csv_dumper_890 = new("./depth890.csv");
    cstatus_csv_dumper_890 = new("./chan_status890.csv");
    fifo_monitor_890 = new(fifo_csv_dumper_890,fifo_intf_890,cstatus_csv_dumper_890);
    fifo_csv_dumper_891 = new("./depth891.csv");
    cstatus_csv_dumper_891 = new("./chan_status891.csv");
    fifo_monitor_891 = new(fifo_csv_dumper_891,fifo_intf_891,cstatus_csv_dumper_891);
    fifo_csv_dumper_892 = new("./depth892.csv");
    cstatus_csv_dumper_892 = new("./chan_status892.csv");
    fifo_monitor_892 = new(fifo_csv_dumper_892,fifo_intf_892,cstatus_csv_dumper_892);
    fifo_csv_dumper_893 = new("./depth893.csv");
    cstatus_csv_dumper_893 = new("./chan_status893.csv");
    fifo_monitor_893 = new(fifo_csv_dumper_893,fifo_intf_893,cstatus_csv_dumper_893);
    fifo_csv_dumper_894 = new("./depth894.csv");
    cstatus_csv_dumper_894 = new("./chan_status894.csv");
    fifo_monitor_894 = new(fifo_csv_dumper_894,fifo_intf_894,cstatus_csv_dumper_894);
    fifo_csv_dumper_895 = new("./depth895.csv");
    cstatus_csv_dumper_895 = new("./chan_status895.csv");
    fifo_monitor_895 = new(fifo_csv_dumper_895,fifo_intf_895,cstatus_csv_dumper_895);
    fifo_csv_dumper_896 = new("./depth896.csv");
    cstatus_csv_dumper_896 = new("./chan_status896.csv");
    fifo_monitor_896 = new(fifo_csv_dumper_896,fifo_intf_896,cstatus_csv_dumper_896);
    fifo_csv_dumper_897 = new("./depth897.csv");
    cstatus_csv_dumper_897 = new("./chan_status897.csv");
    fifo_monitor_897 = new(fifo_csv_dumper_897,fifo_intf_897,cstatus_csv_dumper_897);
    fifo_csv_dumper_898 = new("./depth898.csv");
    cstatus_csv_dumper_898 = new("./chan_status898.csv");
    fifo_monitor_898 = new(fifo_csv_dumper_898,fifo_intf_898,cstatus_csv_dumper_898);
    fifo_csv_dumper_899 = new("./depth899.csv");
    cstatus_csv_dumper_899 = new("./chan_status899.csv");
    fifo_monitor_899 = new(fifo_csv_dumper_899,fifo_intf_899,cstatus_csv_dumper_899);
    fifo_csv_dumper_900 = new("./depth900.csv");
    cstatus_csv_dumper_900 = new("./chan_status900.csv");
    fifo_monitor_900 = new(fifo_csv_dumper_900,fifo_intf_900,cstatus_csv_dumper_900);
    fifo_csv_dumper_901 = new("./depth901.csv");
    cstatus_csv_dumper_901 = new("./chan_status901.csv");
    fifo_monitor_901 = new(fifo_csv_dumper_901,fifo_intf_901,cstatus_csv_dumper_901);
    fifo_csv_dumper_902 = new("./depth902.csv");
    cstatus_csv_dumper_902 = new("./chan_status902.csv");
    fifo_monitor_902 = new(fifo_csv_dumper_902,fifo_intf_902,cstatus_csv_dumper_902);
    fifo_csv_dumper_903 = new("./depth903.csv");
    cstatus_csv_dumper_903 = new("./chan_status903.csv");
    fifo_monitor_903 = new(fifo_csv_dumper_903,fifo_intf_903,cstatus_csv_dumper_903);
    fifo_csv_dumper_904 = new("./depth904.csv");
    cstatus_csv_dumper_904 = new("./chan_status904.csv");
    fifo_monitor_904 = new(fifo_csv_dumper_904,fifo_intf_904,cstatus_csv_dumper_904);
    fifo_csv_dumper_905 = new("./depth905.csv");
    cstatus_csv_dumper_905 = new("./chan_status905.csv");
    fifo_monitor_905 = new(fifo_csv_dumper_905,fifo_intf_905,cstatus_csv_dumper_905);
    fifo_csv_dumper_906 = new("./depth906.csv");
    cstatus_csv_dumper_906 = new("./chan_status906.csv");
    fifo_monitor_906 = new(fifo_csv_dumper_906,fifo_intf_906,cstatus_csv_dumper_906);
    fifo_csv_dumper_907 = new("./depth907.csv");
    cstatus_csv_dumper_907 = new("./chan_status907.csv");
    fifo_monitor_907 = new(fifo_csv_dumper_907,fifo_intf_907,cstatus_csv_dumper_907);
    fifo_csv_dumper_908 = new("./depth908.csv");
    cstatus_csv_dumper_908 = new("./chan_status908.csv");
    fifo_monitor_908 = new(fifo_csv_dumper_908,fifo_intf_908,cstatus_csv_dumper_908);
    fifo_csv_dumper_909 = new("./depth909.csv");
    cstatus_csv_dumper_909 = new("./chan_status909.csv");
    fifo_monitor_909 = new(fifo_csv_dumper_909,fifo_intf_909,cstatus_csv_dumper_909);
    fifo_csv_dumper_910 = new("./depth910.csv");
    cstatus_csv_dumper_910 = new("./chan_status910.csv");
    fifo_monitor_910 = new(fifo_csv_dumper_910,fifo_intf_910,cstatus_csv_dumper_910);
    fifo_csv_dumper_911 = new("./depth911.csv");
    cstatus_csv_dumper_911 = new("./chan_status911.csv");
    fifo_monitor_911 = new(fifo_csv_dumper_911,fifo_intf_911,cstatus_csv_dumper_911);
    fifo_csv_dumper_912 = new("./depth912.csv");
    cstatus_csv_dumper_912 = new("./chan_status912.csv");
    fifo_monitor_912 = new(fifo_csv_dumper_912,fifo_intf_912,cstatus_csv_dumper_912);
    fifo_csv_dumper_913 = new("./depth913.csv");
    cstatus_csv_dumper_913 = new("./chan_status913.csv");
    fifo_monitor_913 = new(fifo_csv_dumper_913,fifo_intf_913,cstatus_csv_dumper_913);
    fifo_csv_dumper_914 = new("./depth914.csv");
    cstatus_csv_dumper_914 = new("./chan_status914.csv");
    fifo_monitor_914 = new(fifo_csv_dumper_914,fifo_intf_914,cstatus_csv_dumper_914);
    fifo_csv_dumper_915 = new("./depth915.csv");
    cstatus_csv_dumper_915 = new("./chan_status915.csv");
    fifo_monitor_915 = new(fifo_csv_dumper_915,fifo_intf_915,cstatus_csv_dumper_915);
    fifo_csv_dumper_916 = new("./depth916.csv");
    cstatus_csv_dumper_916 = new("./chan_status916.csv");
    fifo_monitor_916 = new(fifo_csv_dumper_916,fifo_intf_916,cstatus_csv_dumper_916);
    fifo_csv_dumper_917 = new("./depth917.csv");
    cstatus_csv_dumper_917 = new("./chan_status917.csv");
    fifo_monitor_917 = new(fifo_csv_dumper_917,fifo_intf_917,cstatus_csv_dumper_917);
    fifo_csv_dumper_918 = new("./depth918.csv");
    cstatus_csv_dumper_918 = new("./chan_status918.csv");
    fifo_monitor_918 = new(fifo_csv_dumper_918,fifo_intf_918,cstatus_csv_dumper_918);
    fifo_csv_dumper_919 = new("./depth919.csv");
    cstatus_csv_dumper_919 = new("./chan_status919.csv");
    fifo_monitor_919 = new(fifo_csv_dumper_919,fifo_intf_919,cstatus_csv_dumper_919);
    fifo_csv_dumper_920 = new("./depth920.csv");
    cstatus_csv_dumper_920 = new("./chan_status920.csv");
    fifo_monitor_920 = new(fifo_csv_dumper_920,fifo_intf_920,cstatus_csv_dumper_920);
    fifo_csv_dumper_921 = new("./depth921.csv");
    cstatus_csv_dumper_921 = new("./chan_status921.csv");
    fifo_monitor_921 = new(fifo_csv_dumper_921,fifo_intf_921,cstatus_csv_dumper_921);
    fifo_csv_dumper_922 = new("./depth922.csv");
    cstatus_csv_dumper_922 = new("./chan_status922.csv");
    fifo_monitor_922 = new(fifo_csv_dumper_922,fifo_intf_922,cstatus_csv_dumper_922);
    fifo_csv_dumper_923 = new("./depth923.csv");
    cstatus_csv_dumper_923 = new("./chan_status923.csv");
    fifo_monitor_923 = new(fifo_csv_dumper_923,fifo_intf_923,cstatus_csv_dumper_923);
    fifo_csv_dumper_924 = new("./depth924.csv");
    cstatus_csv_dumper_924 = new("./chan_status924.csv");
    fifo_monitor_924 = new(fifo_csv_dumper_924,fifo_intf_924,cstatus_csv_dumper_924);
    fifo_csv_dumper_925 = new("./depth925.csv");
    cstatus_csv_dumper_925 = new("./chan_status925.csv");
    fifo_monitor_925 = new(fifo_csv_dumper_925,fifo_intf_925,cstatus_csv_dumper_925);
    fifo_csv_dumper_926 = new("./depth926.csv");
    cstatus_csv_dumper_926 = new("./chan_status926.csv");
    fifo_monitor_926 = new(fifo_csv_dumper_926,fifo_intf_926,cstatus_csv_dumper_926);
    fifo_csv_dumper_927 = new("./depth927.csv");
    cstatus_csv_dumper_927 = new("./chan_status927.csv");
    fifo_monitor_927 = new(fifo_csv_dumper_927,fifo_intf_927,cstatus_csv_dumper_927);
    fifo_csv_dumper_928 = new("./depth928.csv");
    cstatus_csv_dumper_928 = new("./chan_status928.csv");
    fifo_monitor_928 = new(fifo_csv_dumper_928,fifo_intf_928,cstatus_csv_dumper_928);
    fifo_csv_dumper_929 = new("./depth929.csv");
    cstatus_csv_dumper_929 = new("./chan_status929.csv");
    fifo_monitor_929 = new(fifo_csv_dumper_929,fifo_intf_929,cstatus_csv_dumper_929);
    fifo_csv_dumper_930 = new("./depth930.csv");
    cstatus_csv_dumper_930 = new("./chan_status930.csv");
    fifo_monitor_930 = new(fifo_csv_dumper_930,fifo_intf_930,cstatus_csv_dumper_930);
    fifo_csv_dumper_931 = new("./depth931.csv");
    cstatus_csv_dumper_931 = new("./chan_status931.csv");
    fifo_monitor_931 = new(fifo_csv_dumper_931,fifo_intf_931,cstatus_csv_dumper_931);
    fifo_csv_dumper_932 = new("./depth932.csv");
    cstatus_csv_dumper_932 = new("./chan_status932.csv");
    fifo_monitor_932 = new(fifo_csv_dumper_932,fifo_intf_932,cstatus_csv_dumper_932);
    fifo_csv_dumper_933 = new("./depth933.csv");
    cstatus_csv_dumper_933 = new("./chan_status933.csv");
    fifo_monitor_933 = new(fifo_csv_dumper_933,fifo_intf_933,cstatus_csv_dumper_933);
    fifo_csv_dumper_934 = new("./depth934.csv");
    cstatus_csv_dumper_934 = new("./chan_status934.csv");
    fifo_monitor_934 = new(fifo_csv_dumper_934,fifo_intf_934,cstatus_csv_dumper_934);
    fifo_csv_dumper_935 = new("./depth935.csv");
    cstatus_csv_dumper_935 = new("./chan_status935.csv");
    fifo_monitor_935 = new(fifo_csv_dumper_935,fifo_intf_935,cstatus_csv_dumper_935);
    fifo_csv_dumper_936 = new("./depth936.csv");
    cstatus_csv_dumper_936 = new("./chan_status936.csv");
    fifo_monitor_936 = new(fifo_csv_dumper_936,fifo_intf_936,cstatus_csv_dumper_936);
    fifo_csv_dumper_937 = new("./depth937.csv");
    cstatus_csv_dumper_937 = new("./chan_status937.csv");
    fifo_monitor_937 = new(fifo_csv_dumper_937,fifo_intf_937,cstatus_csv_dumper_937);
    fifo_csv_dumper_938 = new("./depth938.csv");
    cstatus_csv_dumper_938 = new("./chan_status938.csv");
    fifo_monitor_938 = new(fifo_csv_dumper_938,fifo_intf_938,cstatus_csv_dumper_938);
    fifo_csv_dumper_939 = new("./depth939.csv");
    cstatus_csv_dumper_939 = new("./chan_status939.csv");
    fifo_monitor_939 = new(fifo_csv_dumper_939,fifo_intf_939,cstatus_csv_dumper_939);
    fifo_csv_dumper_940 = new("./depth940.csv");
    cstatus_csv_dumper_940 = new("./chan_status940.csv");
    fifo_monitor_940 = new(fifo_csv_dumper_940,fifo_intf_940,cstatus_csv_dumper_940);
    fifo_csv_dumper_941 = new("./depth941.csv");
    cstatus_csv_dumper_941 = new("./chan_status941.csv");
    fifo_monitor_941 = new(fifo_csv_dumper_941,fifo_intf_941,cstatus_csv_dumper_941);
    fifo_csv_dumper_942 = new("./depth942.csv");
    cstatus_csv_dumper_942 = new("./chan_status942.csv");
    fifo_monitor_942 = new(fifo_csv_dumper_942,fifo_intf_942,cstatus_csv_dumper_942);
    fifo_csv_dumper_943 = new("./depth943.csv");
    cstatus_csv_dumper_943 = new("./chan_status943.csv");
    fifo_monitor_943 = new(fifo_csv_dumper_943,fifo_intf_943,cstatus_csv_dumper_943);
    fifo_csv_dumper_944 = new("./depth944.csv");
    cstatus_csv_dumper_944 = new("./chan_status944.csv");
    fifo_monitor_944 = new(fifo_csv_dumper_944,fifo_intf_944,cstatus_csv_dumper_944);
    fifo_csv_dumper_945 = new("./depth945.csv");
    cstatus_csv_dumper_945 = new("./chan_status945.csv");
    fifo_monitor_945 = new(fifo_csv_dumper_945,fifo_intf_945,cstatus_csv_dumper_945);
    fifo_csv_dumper_946 = new("./depth946.csv");
    cstatus_csv_dumper_946 = new("./chan_status946.csv");
    fifo_monitor_946 = new(fifo_csv_dumper_946,fifo_intf_946,cstatus_csv_dumper_946);
    fifo_csv_dumper_947 = new("./depth947.csv");
    cstatus_csv_dumper_947 = new("./chan_status947.csv");
    fifo_monitor_947 = new(fifo_csv_dumper_947,fifo_intf_947,cstatus_csv_dumper_947);
    fifo_csv_dumper_948 = new("./depth948.csv");
    cstatus_csv_dumper_948 = new("./chan_status948.csv");
    fifo_monitor_948 = new(fifo_csv_dumper_948,fifo_intf_948,cstatus_csv_dumper_948);
    fifo_csv_dumper_949 = new("./depth949.csv");
    cstatus_csv_dumper_949 = new("./chan_status949.csv");
    fifo_monitor_949 = new(fifo_csv_dumper_949,fifo_intf_949,cstatus_csv_dumper_949);
    fifo_csv_dumper_950 = new("./depth950.csv");
    cstatus_csv_dumper_950 = new("./chan_status950.csv");
    fifo_monitor_950 = new(fifo_csv_dumper_950,fifo_intf_950,cstatus_csv_dumper_950);
    fifo_csv_dumper_951 = new("./depth951.csv");
    cstatus_csv_dumper_951 = new("./chan_status951.csv");
    fifo_monitor_951 = new(fifo_csv_dumper_951,fifo_intf_951,cstatus_csv_dumper_951);
    fifo_csv_dumper_952 = new("./depth952.csv");
    cstatus_csv_dumper_952 = new("./chan_status952.csv");
    fifo_monitor_952 = new(fifo_csv_dumper_952,fifo_intf_952,cstatus_csv_dumper_952);
    fifo_csv_dumper_953 = new("./depth953.csv");
    cstatus_csv_dumper_953 = new("./chan_status953.csv");
    fifo_monitor_953 = new(fifo_csv_dumper_953,fifo_intf_953,cstatus_csv_dumper_953);
    fifo_csv_dumper_954 = new("./depth954.csv");
    cstatus_csv_dumper_954 = new("./chan_status954.csv");
    fifo_monitor_954 = new(fifo_csv_dumper_954,fifo_intf_954,cstatus_csv_dumper_954);
    fifo_csv_dumper_955 = new("./depth955.csv");
    cstatus_csv_dumper_955 = new("./chan_status955.csv");
    fifo_monitor_955 = new(fifo_csv_dumper_955,fifo_intf_955,cstatus_csv_dumper_955);
    fifo_csv_dumper_956 = new("./depth956.csv");
    cstatus_csv_dumper_956 = new("./chan_status956.csv");
    fifo_monitor_956 = new(fifo_csv_dumper_956,fifo_intf_956,cstatus_csv_dumper_956);
    fifo_csv_dumper_957 = new("./depth957.csv");
    cstatus_csv_dumper_957 = new("./chan_status957.csv");
    fifo_monitor_957 = new(fifo_csv_dumper_957,fifo_intf_957,cstatus_csv_dumper_957);
    fifo_csv_dumper_958 = new("./depth958.csv");
    cstatus_csv_dumper_958 = new("./chan_status958.csv");
    fifo_monitor_958 = new(fifo_csv_dumper_958,fifo_intf_958,cstatus_csv_dumper_958);
    fifo_csv_dumper_959 = new("./depth959.csv");
    cstatus_csv_dumper_959 = new("./chan_status959.csv");
    fifo_monitor_959 = new(fifo_csv_dumper_959,fifo_intf_959,cstatus_csv_dumper_959);
    fifo_csv_dumper_960 = new("./depth960.csv");
    cstatus_csv_dumper_960 = new("./chan_status960.csv");
    fifo_monitor_960 = new(fifo_csv_dumper_960,fifo_intf_960,cstatus_csv_dumper_960);
    fifo_csv_dumper_961 = new("./depth961.csv");
    cstatus_csv_dumper_961 = new("./chan_status961.csv");
    fifo_monitor_961 = new(fifo_csv_dumper_961,fifo_intf_961,cstatus_csv_dumper_961);
    fifo_csv_dumper_962 = new("./depth962.csv");
    cstatus_csv_dumper_962 = new("./chan_status962.csv");
    fifo_monitor_962 = new(fifo_csv_dumper_962,fifo_intf_962,cstatus_csv_dumper_962);
    fifo_csv_dumper_963 = new("./depth963.csv");
    cstatus_csv_dumper_963 = new("./chan_status963.csv");
    fifo_monitor_963 = new(fifo_csv_dumper_963,fifo_intf_963,cstatus_csv_dumper_963);
    fifo_csv_dumper_964 = new("./depth964.csv");
    cstatus_csv_dumper_964 = new("./chan_status964.csv");
    fifo_monitor_964 = new(fifo_csv_dumper_964,fifo_intf_964,cstatus_csv_dumper_964);
    fifo_csv_dumper_965 = new("./depth965.csv");
    cstatus_csv_dumper_965 = new("./chan_status965.csv");
    fifo_monitor_965 = new(fifo_csv_dumper_965,fifo_intf_965,cstatus_csv_dumper_965);
    fifo_csv_dumper_966 = new("./depth966.csv");
    cstatus_csv_dumper_966 = new("./chan_status966.csv");
    fifo_monitor_966 = new(fifo_csv_dumper_966,fifo_intf_966,cstatus_csv_dumper_966);
    fifo_csv_dumper_967 = new("./depth967.csv");
    cstatus_csv_dumper_967 = new("./chan_status967.csv");
    fifo_monitor_967 = new(fifo_csv_dumper_967,fifo_intf_967,cstatus_csv_dumper_967);
    fifo_csv_dumper_968 = new("./depth968.csv");
    cstatus_csv_dumper_968 = new("./chan_status968.csv");
    fifo_monitor_968 = new(fifo_csv_dumper_968,fifo_intf_968,cstatus_csv_dumper_968);
    fifo_csv_dumper_969 = new("./depth969.csv");
    cstatus_csv_dumper_969 = new("./chan_status969.csv");
    fifo_monitor_969 = new(fifo_csv_dumper_969,fifo_intf_969,cstatus_csv_dumper_969);
    fifo_csv_dumper_970 = new("./depth970.csv");
    cstatus_csv_dumper_970 = new("./chan_status970.csv");
    fifo_monitor_970 = new(fifo_csv_dumper_970,fifo_intf_970,cstatus_csv_dumper_970);
    fifo_csv_dumper_971 = new("./depth971.csv");
    cstatus_csv_dumper_971 = new("./chan_status971.csv");
    fifo_monitor_971 = new(fifo_csv_dumper_971,fifo_intf_971,cstatus_csv_dumper_971);
    fifo_csv_dumper_972 = new("./depth972.csv");
    cstatus_csv_dumper_972 = new("./chan_status972.csv");
    fifo_monitor_972 = new(fifo_csv_dumper_972,fifo_intf_972,cstatus_csv_dumper_972);
    fifo_csv_dumper_973 = new("./depth973.csv");
    cstatus_csv_dumper_973 = new("./chan_status973.csv");
    fifo_monitor_973 = new(fifo_csv_dumper_973,fifo_intf_973,cstatus_csv_dumper_973);
    fifo_csv_dumper_974 = new("./depth974.csv");
    cstatus_csv_dumper_974 = new("./chan_status974.csv");
    fifo_monitor_974 = new(fifo_csv_dumper_974,fifo_intf_974,cstatus_csv_dumper_974);
    fifo_csv_dumper_975 = new("./depth975.csv");
    cstatus_csv_dumper_975 = new("./chan_status975.csv");
    fifo_monitor_975 = new(fifo_csv_dumper_975,fifo_intf_975,cstatus_csv_dumper_975);
    fifo_csv_dumper_976 = new("./depth976.csv");
    cstatus_csv_dumper_976 = new("./chan_status976.csv");
    fifo_monitor_976 = new(fifo_csv_dumper_976,fifo_intf_976,cstatus_csv_dumper_976);
    fifo_csv_dumper_977 = new("./depth977.csv");
    cstatus_csv_dumper_977 = new("./chan_status977.csv");
    fifo_monitor_977 = new(fifo_csv_dumper_977,fifo_intf_977,cstatus_csv_dumper_977);
    fifo_csv_dumper_978 = new("./depth978.csv");
    cstatus_csv_dumper_978 = new("./chan_status978.csv");
    fifo_monitor_978 = new(fifo_csv_dumper_978,fifo_intf_978,cstatus_csv_dumper_978);
    fifo_csv_dumper_979 = new("./depth979.csv");
    cstatus_csv_dumper_979 = new("./chan_status979.csv");
    fifo_monitor_979 = new(fifo_csv_dumper_979,fifo_intf_979,cstatus_csv_dumper_979);
    fifo_csv_dumper_980 = new("./depth980.csv");
    cstatus_csv_dumper_980 = new("./chan_status980.csv");
    fifo_monitor_980 = new(fifo_csv_dumper_980,fifo_intf_980,cstatus_csv_dumper_980);
    fifo_csv_dumper_981 = new("./depth981.csv");
    cstatus_csv_dumper_981 = new("./chan_status981.csv");
    fifo_monitor_981 = new(fifo_csv_dumper_981,fifo_intf_981,cstatus_csv_dumper_981);
    fifo_csv_dumper_982 = new("./depth982.csv");
    cstatus_csv_dumper_982 = new("./chan_status982.csv");
    fifo_monitor_982 = new(fifo_csv_dumper_982,fifo_intf_982,cstatus_csv_dumper_982);
    fifo_csv_dumper_983 = new("./depth983.csv");
    cstatus_csv_dumper_983 = new("./chan_status983.csv");
    fifo_monitor_983 = new(fifo_csv_dumper_983,fifo_intf_983,cstatus_csv_dumper_983);
    fifo_csv_dumper_984 = new("./depth984.csv");
    cstatus_csv_dumper_984 = new("./chan_status984.csv");
    fifo_monitor_984 = new(fifo_csv_dumper_984,fifo_intf_984,cstatus_csv_dumper_984);
    fifo_csv_dumper_985 = new("./depth985.csv");
    cstatus_csv_dumper_985 = new("./chan_status985.csv");
    fifo_monitor_985 = new(fifo_csv_dumper_985,fifo_intf_985,cstatus_csv_dumper_985);
    fifo_csv_dumper_986 = new("./depth986.csv");
    cstatus_csv_dumper_986 = new("./chan_status986.csv");
    fifo_monitor_986 = new(fifo_csv_dumper_986,fifo_intf_986,cstatus_csv_dumper_986);
    fifo_csv_dumper_987 = new("./depth987.csv");
    cstatus_csv_dumper_987 = new("./chan_status987.csv");
    fifo_monitor_987 = new(fifo_csv_dumper_987,fifo_intf_987,cstatus_csv_dumper_987);
    fifo_csv_dumper_988 = new("./depth988.csv");
    cstatus_csv_dumper_988 = new("./chan_status988.csv");
    fifo_monitor_988 = new(fifo_csv_dumper_988,fifo_intf_988,cstatus_csv_dumper_988);
    fifo_csv_dumper_989 = new("./depth989.csv");
    cstatus_csv_dumper_989 = new("./chan_status989.csv");
    fifo_monitor_989 = new(fifo_csv_dumper_989,fifo_intf_989,cstatus_csv_dumper_989);
    fifo_csv_dumper_990 = new("./depth990.csv");
    cstatus_csv_dumper_990 = new("./chan_status990.csv");
    fifo_monitor_990 = new(fifo_csv_dumper_990,fifo_intf_990,cstatus_csv_dumper_990);
    fifo_csv_dumper_991 = new("./depth991.csv");
    cstatus_csv_dumper_991 = new("./chan_status991.csv");
    fifo_monitor_991 = new(fifo_csv_dumper_991,fifo_intf_991,cstatus_csv_dumper_991);
    fifo_csv_dumper_992 = new("./depth992.csv");
    cstatus_csv_dumper_992 = new("./chan_status992.csv");
    fifo_monitor_992 = new(fifo_csv_dumper_992,fifo_intf_992,cstatus_csv_dumper_992);
    fifo_csv_dumper_993 = new("./depth993.csv");
    cstatus_csv_dumper_993 = new("./chan_status993.csv");
    fifo_monitor_993 = new(fifo_csv_dumper_993,fifo_intf_993,cstatus_csv_dumper_993);
    fifo_csv_dumper_994 = new("./depth994.csv");
    cstatus_csv_dumper_994 = new("./chan_status994.csv");
    fifo_monitor_994 = new(fifo_csv_dumper_994,fifo_intf_994,cstatus_csv_dumper_994);
    fifo_csv_dumper_995 = new("./depth995.csv");
    cstatus_csv_dumper_995 = new("./chan_status995.csv");
    fifo_monitor_995 = new(fifo_csv_dumper_995,fifo_intf_995,cstatus_csv_dumper_995);
    fifo_csv_dumper_996 = new("./depth996.csv");
    cstatus_csv_dumper_996 = new("./chan_status996.csv");
    fifo_monitor_996 = new(fifo_csv_dumper_996,fifo_intf_996,cstatus_csv_dumper_996);
    fifo_csv_dumper_997 = new("./depth997.csv");
    cstatus_csv_dumper_997 = new("./chan_status997.csv");
    fifo_monitor_997 = new(fifo_csv_dumper_997,fifo_intf_997,cstatus_csv_dumper_997);
    fifo_csv_dumper_998 = new("./depth998.csv");
    cstatus_csv_dumper_998 = new("./chan_status998.csv");
    fifo_monitor_998 = new(fifo_csv_dumper_998,fifo_intf_998,cstatus_csv_dumper_998);
    fifo_csv_dumper_999 = new("./depth999.csv");
    cstatus_csv_dumper_999 = new("./chan_status999.csv");
    fifo_monitor_999 = new(fifo_csv_dumper_999,fifo_intf_999,cstatus_csv_dumper_999);
    fifo_csv_dumper_1000 = new("./depth1000.csv");
    cstatus_csv_dumper_1000 = new("./chan_status1000.csv");
    fifo_monitor_1000 = new(fifo_csv_dumper_1000,fifo_intf_1000,cstatus_csv_dumper_1000);
    fifo_csv_dumper_1001 = new("./depth1001.csv");
    cstatus_csv_dumper_1001 = new("./chan_status1001.csv");
    fifo_monitor_1001 = new(fifo_csv_dumper_1001,fifo_intf_1001,cstatus_csv_dumper_1001);
    fifo_csv_dumper_1002 = new("./depth1002.csv");
    cstatus_csv_dumper_1002 = new("./chan_status1002.csv");
    fifo_monitor_1002 = new(fifo_csv_dumper_1002,fifo_intf_1002,cstatus_csv_dumper_1002);
    fifo_csv_dumper_1003 = new("./depth1003.csv");
    cstatus_csv_dumper_1003 = new("./chan_status1003.csv");
    fifo_monitor_1003 = new(fifo_csv_dumper_1003,fifo_intf_1003,cstatus_csv_dumper_1003);
    fifo_csv_dumper_1004 = new("./depth1004.csv");
    cstatus_csv_dumper_1004 = new("./chan_status1004.csv");
    fifo_monitor_1004 = new(fifo_csv_dumper_1004,fifo_intf_1004,cstatus_csv_dumper_1004);
    fifo_csv_dumper_1005 = new("./depth1005.csv");
    cstatus_csv_dumper_1005 = new("./chan_status1005.csv");
    fifo_monitor_1005 = new(fifo_csv_dumper_1005,fifo_intf_1005,cstatus_csv_dumper_1005);
    fifo_csv_dumper_1006 = new("./depth1006.csv");
    cstatus_csv_dumper_1006 = new("./chan_status1006.csv");
    fifo_monitor_1006 = new(fifo_csv_dumper_1006,fifo_intf_1006,cstatus_csv_dumper_1006);
    fifo_csv_dumper_1007 = new("./depth1007.csv");
    cstatus_csv_dumper_1007 = new("./chan_status1007.csv");
    fifo_monitor_1007 = new(fifo_csv_dumper_1007,fifo_intf_1007,cstatus_csv_dumper_1007);
    fifo_csv_dumper_1008 = new("./depth1008.csv");
    cstatus_csv_dumper_1008 = new("./chan_status1008.csv");
    fifo_monitor_1008 = new(fifo_csv_dumper_1008,fifo_intf_1008,cstatus_csv_dumper_1008);
    fifo_csv_dumper_1009 = new("./depth1009.csv");
    cstatus_csv_dumper_1009 = new("./chan_status1009.csv");
    fifo_monitor_1009 = new(fifo_csv_dumper_1009,fifo_intf_1009,cstatus_csv_dumper_1009);
    fifo_csv_dumper_1010 = new("./depth1010.csv");
    cstatus_csv_dumper_1010 = new("./chan_status1010.csv");
    fifo_monitor_1010 = new(fifo_csv_dumper_1010,fifo_intf_1010,cstatus_csv_dumper_1010);
    fifo_csv_dumper_1011 = new("./depth1011.csv");
    cstatus_csv_dumper_1011 = new("./chan_status1011.csv");
    fifo_monitor_1011 = new(fifo_csv_dumper_1011,fifo_intf_1011,cstatus_csv_dumper_1011);
    fifo_csv_dumper_1012 = new("./depth1012.csv");
    cstatus_csv_dumper_1012 = new("./chan_status1012.csv");
    fifo_monitor_1012 = new(fifo_csv_dumper_1012,fifo_intf_1012,cstatus_csv_dumper_1012);
    fifo_csv_dumper_1013 = new("./depth1013.csv");
    cstatus_csv_dumper_1013 = new("./chan_status1013.csv");
    fifo_monitor_1013 = new(fifo_csv_dumper_1013,fifo_intf_1013,cstatus_csv_dumper_1013);
    fifo_csv_dumper_1014 = new("./depth1014.csv");
    cstatus_csv_dumper_1014 = new("./chan_status1014.csv");
    fifo_monitor_1014 = new(fifo_csv_dumper_1014,fifo_intf_1014,cstatus_csv_dumper_1014);
    fifo_csv_dumper_1015 = new("./depth1015.csv");
    cstatus_csv_dumper_1015 = new("./chan_status1015.csv");
    fifo_monitor_1015 = new(fifo_csv_dumper_1015,fifo_intf_1015,cstatus_csv_dumper_1015);
    fifo_csv_dumper_1016 = new("./depth1016.csv");
    cstatus_csv_dumper_1016 = new("./chan_status1016.csv");
    fifo_monitor_1016 = new(fifo_csv_dumper_1016,fifo_intf_1016,cstatus_csv_dumper_1016);
    fifo_csv_dumper_1017 = new("./depth1017.csv");
    cstatus_csv_dumper_1017 = new("./chan_status1017.csv");
    fifo_monitor_1017 = new(fifo_csv_dumper_1017,fifo_intf_1017,cstatus_csv_dumper_1017);
    fifo_csv_dumper_1018 = new("./depth1018.csv");
    cstatus_csv_dumper_1018 = new("./chan_status1018.csv");
    fifo_monitor_1018 = new(fifo_csv_dumper_1018,fifo_intf_1018,cstatus_csv_dumper_1018);
    fifo_csv_dumper_1019 = new("./depth1019.csv");
    cstatus_csv_dumper_1019 = new("./chan_status1019.csv");
    fifo_monitor_1019 = new(fifo_csv_dumper_1019,fifo_intf_1019,cstatus_csv_dumper_1019);
    fifo_csv_dumper_1020 = new("./depth1020.csv");
    cstatus_csv_dumper_1020 = new("./chan_status1020.csv");
    fifo_monitor_1020 = new(fifo_csv_dumper_1020,fifo_intf_1020,cstatus_csv_dumper_1020);
    fifo_csv_dumper_1021 = new("./depth1021.csv");
    cstatus_csv_dumper_1021 = new("./chan_status1021.csv");
    fifo_monitor_1021 = new(fifo_csv_dumper_1021,fifo_intf_1021,cstatus_csv_dumper_1021);
    fifo_csv_dumper_1022 = new("./depth1022.csv");
    cstatus_csv_dumper_1022 = new("./chan_status1022.csv");
    fifo_monitor_1022 = new(fifo_csv_dumper_1022,fifo_intf_1022,cstatus_csv_dumper_1022);
    fifo_csv_dumper_1023 = new("./depth1023.csv");
    cstatus_csv_dumper_1023 = new("./chan_status1023.csv");
    fifo_monitor_1023 = new(fifo_csv_dumper_1023,fifo_intf_1023,cstatus_csv_dumper_1023);
    fifo_csv_dumper_1024 = new("./depth1024.csv");
    cstatus_csv_dumper_1024 = new("./chan_status1024.csv");
    fifo_monitor_1024 = new(fifo_csv_dumper_1024,fifo_intf_1024,cstatus_csv_dumper_1024);
    fifo_csv_dumper_1025 = new("./depth1025.csv");
    cstatus_csv_dumper_1025 = new("./chan_status1025.csv");
    fifo_monitor_1025 = new(fifo_csv_dumper_1025,fifo_intf_1025,cstatus_csv_dumper_1025);
    fifo_csv_dumper_1026 = new("./depth1026.csv");
    cstatus_csv_dumper_1026 = new("./chan_status1026.csv");
    fifo_monitor_1026 = new(fifo_csv_dumper_1026,fifo_intf_1026,cstatus_csv_dumper_1026);
    fifo_csv_dumper_1027 = new("./depth1027.csv");
    cstatus_csv_dumper_1027 = new("./chan_status1027.csv");
    fifo_monitor_1027 = new(fifo_csv_dumper_1027,fifo_intf_1027,cstatus_csv_dumper_1027);
    fifo_csv_dumper_1028 = new("./depth1028.csv");
    cstatus_csv_dumper_1028 = new("./chan_status1028.csv");
    fifo_monitor_1028 = new(fifo_csv_dumper_1028,fifo_intf_1028,cstatus_csv_dumper_1028);
    fifo_csv_dumper_1029 = new("./depth1029.csv");
    cstatus_csv_dumper_1029 = new("./chan_status1029.csv");
    fifo_monitor_1029 = new(fifo_csv_dumper_1029,fifo_intf_1029,cstatus_csv_dumper_1029);
    fifo_csv_dumper_1030 = new("./depth1030.csv");
    cstatus_csv_dumper_1030 = new("./chan_status1030.csv");
    fifo_monitor_1030 = new(fifo_csv_dumper_1030,fifo_intf_1030,cstatus_csv_dumper_1030);
    fifo_csv_dumper_1031 = new("./depth1031.csv");
    cstatus_csv_dumper_1031 = new("./chan_status1031.csv");
    fifo_monitor_1031 = new(fifo_csv_dumper_1031,fifo_intf_1031,cstatus_csv_dumper_1031);
    fifo_csv_dumper_1032 = new("./depth1032.csv");
    cstatus_csv_dumper_1032 = new("./chan_status1032.csv");
    fifo_monitor_1032 = new(fifo_csv_dumper_1032,fifo_intf_1032,cstatus_csv_dumper_1032);
    fifo_csv_dumper_1033 = new("./depth1033.csv");
    cstatus_csv_dumper_1033 = new("./chan_status1033.csv");
    fifo_monitor_1033 = new(fifo_csv_dumper_1033,fifo_intf_1033,cstatus_csv_dumper_1033);
    fifo_csv_dumper_1034 = new("./depth1034.csv");
    cstatus_csv_dumper_1034 = new("./chan_status1034.csv");
    fifo_monitor_1034 = new(fifo_csv_dumper_1034,fifo_intf_1034,cstatus_csv_dumper_1034);
    fifo_csv_dumper_1035 = new("./depth1035.csv");
    cstatus_csv_dumper_1035 = new("./chan_status1035.csv");
    fifo_monitor_1035 = new(fifo_csv_dumper_1035,fifo_intf_1035,cstatus_csv_dumper_1035);
    fifo_csv_dumper_1036 = new("./depth1036.csv");
    cstatus_csv_dumper_1036 = new("./chan_status1036.csv");
    fifo_monitor_1036 = new(fifo_csv_dumper_1036,fifo_intf_1036,cstatus_csv_dumper_1036);
    fifo_csv_dumper_1037 = new("./depth1037.csv");
    cstatus_csv_dumper_1037 = new("./chan_status1037.csv");
    fifo_monitor_1037 = new(fifo_csv_dumper_1037,fifo_intf_1037,cstatus_csv_dumper_1037);
    fifo_csv_dumper_1038 = new("./depth1038.csv");
    cstatus_csv_dumper_1038 = new("./chan_status1038.csv");
    fifo_monitor_1038 = new(fifo_csv_dumper_1038,fifo_intf_1038,cstatus_csv_dumper_1038);
    fifo_csv_dumper_1039 = new("./depth1039.csv");
    cstatus_csv_dumper_1039 = new("./chan_status1039.csv");
    fifo_monitor_1039 = new(fifo_csv_dumper_1039,fifo_intf_1039,cstatus_csv_dumper_1039);
    fifo_csv_dumper_1040 = new("./depth1040.csv");
    cstatus_csv_dumper_1040 = new("./chan_status1040.csv");
    fifo_monitor_1040 = new(fifo_csv_dumper_1040,fifo_intf_1040,cstatus_csv_dumper_1040);
    fifo_csv_dumper_1041 = new("./depth1041.csv");
    cstatus_csv_dumper_1041 = new("./chan_status1041.csv");
    fifo_monitor_1041 = new(fifo_csv_dumper_1041,fifo_intf_1041,cstatus_csv_dumper_1041);
    fifo_csv_dumper_1042 = new("./depth1042.csv");
    cstatus_csv_dumper_1042 = new("./chan_status1042.csv");
    fifo_monitor_1042 = new(fifo_csv_dumper_1042,fifo_intf_1042,cstatus_csv_dumper_1042);
    fifo_csv_dumper_1043 = new("./depth1043.csv");
    cstatus_csv_dumper_1043 = new("./chan_status1043.csv");
    fifo_monitor_1043 = new(fifo_csv_dumper_1043,fifo_intf_1043,cstatus_csv_dumper_1043);
    fifo_csv_dumper_1044 = new("./depth1044.csv");
    cstatus_csv_dumper_1044 = new("./chan_status1044.csv");
    fifo_monitor_1044 = new(fifo_csv_dumper_1044,fifo_intf_1044,cstatus_csv_dumper_1044);
    fifo_csv_dumper_1045 = new("./depth1045.csv");
    cstatus_csv_dumper_1045 = new("./chan_status1045.csv");
    fifo_monitor_1045 = new(fifo_csv_dumper_1045,fifo_intf_1045,cstatus_csv_dumper_1045);
    fifo_csv_dumper_1046 = new("./depth1046.csv");
    cstatus_csv_dumper_1046 = new("./chan_status1046.csv");
    fifo_monitor_1046 = new(fifo_csv_dumper_1046,fifo_intf_1046,cstatus_csv_dumper_1046);
    fifo_csv_dumper_1047 = new("./depth1047.csv");
    cstatus_csv_dumper_1047 = new("./chan_status1047.csv");
    fifo_monitor_1047 = new(fifo_csv_dumper_1047,fifo_intf_1047,cstatus_csv_dumper_1047);
    fifo_csv_dumper_1048 = new("./depth1048.csv");
    cstatus_csv_dumper_1048 = new("./chan_status1048.csv");
    fifo_monitor_1048 = new(fifo_csv_dumper_1048,fifo_intf_1048,cstatus_csv_dumper_1048);
    fifo_csv_dumper_1049 = new("./depth1049.csv");
    cstatus_csv_dumper_1049 = new("./chan_status1049.csv");
    fifo_monitor_1049 = new(fifo_csv_dumper_1049,fifo_intf_1049,cstatus_csv_dumper_1049);
    fifo_csv_dumper_1050 = new("./depth1050.csv");
    cstatus_csv_dumper_1050 = new("./chan_status1050.csv");
    fifo_monitor_1050 = new(fifo_csv_dumper_1050,fifo_intf_1050,cstatus_csv_dumper_1050);
    fifo_csv_dumper_1051 = new("./depth1051.csv");
    cstatus_csv_dumper_1051 = new("./chan_status1051.csv");
    fifo_monitor_1051 = new(fifo_csv_dumper_1051,fifo_intf_1051,cstatus_csv_dumper_1051);
    fifo_csv_dumper_1052 = new("./depth1052.csv");
    cstatus_csv_dumper_1052 = new("./chan_status1052.csv");
    fifo_monitor_1052 = new(fifo_csv_dumper_1052,fifo_intf_1052,cstatus_csv_dumper_1052);
    fifo_csv_dumper_1053 = new("./depth1053.csv");
    cstatus_csv_dumper_1053 = new("./chan_status1053.csv");
    fifo_monitor_1053 = new(fifo_csv_dumper_1053,fifo_intf_1053,cstatus_csv_dumper_1053);
    fifo_csv_dumper_1054 = new("./depth1054.csv");
    cstatus_csv_dumper_1054 = new("./chan_status1054.csv");
    fifo_monitor_1054 = new(fifo_csv_dumper_1054,fifo_intf_1054,cstatus_csv_dumper_1054);
    fifo_csv_dumper_1055 = new("./depth1055.csv");
    cstatus_csv_dumper_1055 = new("./chan_status1055.csv");
    fifo_monitor_1055 = new(fifo_csv_dumper_1055,fifo_intf_1055,cstatus_csv_dumper_1055);
    fifo_csv_dumper_1056 = new("./depth1056.csv");
    cstatus_csv_dumper_1056 = new("./chan_status1056.csv");
    fifo_monitor_1056 = new(fifo_csv_dumper_1056,fifo_intf_1056,cstatus_csv_dumper_1056);
    fifo_csv_dumper_1057 = new("./depth1057.csv");
    cstatus_csv_dumper_1057 = new("./chan_status1057.csv");
    fifo_monitor_1057 = new(fifo_csv_dumper_1057,fifo_intf_1057,cstatus_csv_dumper_1057);
    fifo_csv_dumper_1058 = new("./depth1058.csv");
    cstatus_csv_dumper_1058 = new("./chan_status1058.csv");
    fifo_monitor_1058 = new(fifo_csv_dumper_1058,fifo_intf_1058,cstatus_csv_dumper_1058);
    fifo_csv_dumper_1059 = new("./depth1059.csv");
    cstatus_csv_dumper_1059 = new("./chan_status1059.csv");
    fifo_monitor_1059 = new(fifo_csv_dumper_1059,fifo_intf_1059,cstatus_csv_dumper_1059);
    fifo_csv_dumper_1060 = new("./depth1060.csv");
    cstatus_csv_dumper_1060 = new("./chan_status1060.csv");
    fifo_monitor_1060 = new(fifo_csv_dumper_1060,fifo_intf_1060,cstatus_csv_dumper_1060);
    fifo_csv_dumper_1061 = new("./depth1061.csv");
    cstatus_csv_dumper_1061 = new("./chan_status1061.csv");
    fifo_monitor_1061 = new(fifo_csv_dumper_1061,fifo_intf_1061,cstatus_csv_dumper_1061);
    fifo_csv_dumper_1062 = new("./depth1062.csv");
    cstatus_csv_dumper_1062 = new("./chan_status1062.csv");
    fifo_monitor_1062 = new(fifo_csv_dumper_1062,fifo_intf_1062,cstatus_csv_dumper_1062);
    fifo_csv_dumper_1063 = new("./depth1063.csv");
    cstatus_csv_dumper_1063 = new("./chan_status1063.csv");
    fifo_monitor_1063 = new(fifo_csv_dumper_1063,fifo_intf_1063,cstatus_csv_dumper_1063);
    fifo_csv_dumper_1064 = new("./depth1064.csv");
    cstatus_csv_dumper_1064 = new("./chan_status1064.csv");
    fifo_monitor_1064 = new(fifo_csv_dumper_1064,fifo_intf_1064,cstatus_csv_dumper_1064);
    fifo_csv_dumper_1065 = new("./depth1065.csv");
    cstatus_csv_dumper_1065 = new("./chan_status1065.csv");
    fifo_monitor_1065 = new(fifo_csv_dumper_1065,fifo_intf_1065,cstatus_csv_dumper_1065);
    fifo_csv_dumper_1066 = new("./depth1066.csv");
    cstatus_csv_dumper_1066 = new("./chan_status1066.csv");
    fifo_monitor_1066 = new(fifo_csv_dumper_1066,fifo_intf_1066,cstatus_csv_dumper_1066);
    fifo_csv_dumper_1067 = new("./depth1067.csv");
    cstatus_csv_dumper_1067 = new("./chan_status1067.csv");
    fifo_monitor_1067 = new(fifo_csv_dumper_1067,fifo_intf_1067,cstatus_csv_dumper_1067);
    fifo_csv_dumper_1068 = new("./depth1068.csv");
    cstatus_csv_dumper_1068 = new("./chan_status1068.csv");
    fifo_monitor_1068 = new(fifo_csv_dumper_1068,fifo_intf_1068,cstatus_csv_dumper_1068);
    fifo_csv_dumper_1069 = new("./depth1069.csv");
    cstatus_csv_dumper_1069 = new("./chan_status1069.csv");
    fifo_monitor_1069 = new(fifo_csv_dumper_1069,fifo_intf_1069,cstatus_csv_dumper_1069);
    fifo_csv_dumper_1070 = new("./depth1070.csv");
    cstatus_csv_dumper_1070 = new("./chan_status1070.csv");
    fifo_monitor_1070 = new(fifo_csv_dumper_1070,fifo_intf_1070,cstatus_csv_dumper_1070);
    fifo_csv_dumper_1071 = new("./depth1071.csv");
    cstatus_csv_dumper_1071 = new("./chan_status1071.csv");
    fifo_monitor_1071 = new(fifo_csv_dumper_1071,fifo_intf_1071,cstatus_csv_dumper_1071);
    fifo_csv_dumper_1072 = new("./depth1072.csv");
    cstatus_csv_dumper_1072 = new("./chan_status1072.csv");
    fifo_monitor_1072 = new(fifo_csv_dumper_1072,fifo_intf_1072,cstatus_csv_dumper_1072);
    fifo_csv_dumper_1073 = new("./depth1073.csv");
    cstatus_csv_dumper_1073 = new("./chan_status1073.csv");
    fifo_monitor_1073 = new(fifo_csv_dumper_1073,fifo_intf_1073,cstatus_csv_dumper_1073);
    fifo_csv_dumper_1074 = new("./depth1074.csv");
    cstatus_csv_dumper_1074 = new("./chan_status1074.csv");
    fifo_monitor_1074 = new(fifo_csv_dumper_1074,fifo_intf_1074,cstatus_csv_dumper_1074);
    fifo_csv_dumper_1075 = new("./depth1075.csv");
    cstatus_csv_dumper_1075 = new("./chan_status1075.csv");
    fifo_monitor_1075 = new(fifo_csv_dumper_1075,fifo_intf_1075,cstatus_csv_dumper_1075);
    fifo_csv_dumper_1076 = new("./depth1076.csv");
    cstatus_csv_dumper_1076 = new("./chan_status1076.csv");
    fifo_monitor_1076 = new(fifo_csv_dumper_1076,fifo_intf_1076,cstatus_csv_dumper_1076);
    fifo_csv_dumper_1077 = new("./depth1077.csv");
    cstatus_csv_dumper_1077 = new("./chan_status1077.csv");
    fifo_monitor_1077 = new(fifo_csv_dumper_1077,fifo_intf_1077,cstatus_csv_dumper_1077);
    fifo_csv_dumper_1078 = new("./depth1078.csv");
    cstatus_csv_dumper_1078 = new("./chan_status1078.csv");
    fifo_monitor_1078 = new(fifo_csv_dumper_1078,fifo_intf_1078,cstatus_csv_dumper_1078);
    fifo_csv_dumper_1079 = new("./depth1079.csv");
    cstatus_csv_dumper_1079 = new("./chan_status1079.csv");
    fifo_monitor_1079 = new(fifo_csv_dumper_1079,fifo_intf_1079,cstatus_csv_dumper_1079);
    fifo_csv_dumper_1080 = new("./depth1080.csv");
    cstatus_csv_dumper_1080 = new("./chan_status1080.csv");
    fifo_monitor_1080 = new(fifo_csv_dumper_1080,fifo_intf_1080,cstatus_csv_dumper_1080);
    fifo_csv_dumper_1081 = new("./depth1081.csv");
    cstatus_csv_dumper_1081 = new("./chan_status1081.csv");
    fifo_monitor_1081 = new(fifo_csv_dumper_1081,fifo_intf_1081,cstatus_csv_dumper_1081);
    fifo_csv_dumper_1082 = new("./depth1082.csv");
    cstatus_csv_dumper_1082 = new("./chan_status1082.csv");
    fifo_monitor_1082 = new(fifo_csv_dumper_1082,fifo_intf_1082,cstatus_csv_dumper_1082);
    fifo_csv_dumper_1083 = new("./depth1083.csv");
    cstatus_csv_dumper_1083 = new("./chan_status1083.csv");
    fifo_monitor_1083 = new(fifo_csv_dumper_1083,fifo_intf_1083,cstatus_csv_dumper_1083);
    fifo_csv_dumper_1084 = new("./depth1084.csv");
    cstatus_csv_dumper_1084 = new("./chan_status1084.csv");
    fifo_monitor_1084 = new(fifo_csv_dumper_1084,fifo_intf_1084,cstatus_csv_dumper_1084);
    fifo_csv_dumper_1085 = new("./depth1085.csv");
    cstatus_csv_dumper_1085 = new("./chan_status1085.csv");
    fifo_monitor_1085 = new(fifo_csv_dumper_1085,fifo_intf_1085,cstatus_csv_dumper_1085);
    fifo_csv_dumper_1086 = new("./depth1086.csv");
    cstatus_csv_dumper_1086 = new("./chan_status1086.csv");
    fifo_monitor_1086 = new(fifo_csv_dumper_1086,fifo_intf_1086,cstatus_csv_dumper_1086);
    fifo_csv_dumper_1087 = new("./depth1087.csv");
    cstatus_csv_dumper_1087 = new("./chan_status1087.csv");
    fifo_monitor_1087 = new(fifo_csv_dumper_1087,fifo_intf_1087,cstatus_csv_dumper_1087);
    fifo_csv_dumper_1088 = new("./depth1088.csv");
    cstatus_csv_dumper_1088 = new("./chan_status1088.csv");
    fifo_monitor_1088 = new(fifo_csv_dumper_1088,fifo_intf_1088,cstatus_csv_dumper_1088);
    fifo_csv_dumper_1089 = new("./depth1089.csv");
    cstatus_csv_dumper_1089 = new("./chan_status1089.csv");
    fifo_monitor_1089 = new(fifo_csv_dumper_1089,fifo_intf_1089,cstatus_csv_dumper_1089);
    fifo_csv_dumper_1090 = new("./depth1090.csv");
    cstatus_csv_dumper_1090 = new("./chan_status1090.csv");
    fifo_monitor_1090 = new(fifo_csv_dumper_1090,fifo_intf_1090,cstatus_csv_dumper_1090);
    fifo_csv_dumper_1091 = new("./depth1091.csv");
    cstatus_csv_dumper_1091 = new("./chan_status1091.csv");
    fifo_monitor_1091 = new(fifo_csv_dumper_1091,fifo_intf_1091,cstatus_csv_dumper_1091);
    fifo_csv_dumper_1092 = new("./depth1092.csv");
    cstatus_csv_dumper_1092 = new("./chan_status1092.csv");
    fifo_monitor_1092 = new(fifo_csv_dumper_1092,fifo_intf_1092,cstatus_csv_dumper_1092);
    fifo_csv_dumper_1093 = new("./depth1093.csv");
    cstatus_csv_dumper_1093 = new("./chan_status1093.csv");
    fifo_monitor_1093 = new(fifo_csv_dumper_1093,fifo_intf_1093,cstatus_csv_dumper_1093);
    fifo_csv_dumper_1094 = new("./depth1094.csv");
    cstatus_csv_dumper_1094 = new("./chan_status1094.csv");
    fifo_monitor_1094 = new(fifo_csv_dumper_1094,fifo_intf_1094,cstatus_csv_dumper_1094);
    fifo_csv_dumper_1095 = new("./depth1095.csv");
    cstatus_csv_dumper_1095 = new("./chan_status1095.csv");
    fifo_monitor_1095 = new(fifo_csv_dumper_1095,fifo_intf_1095,cstatus_csv_dumper_1095);
    fifo_csv_dumper_1096 = new("./depth1096.csv");
    cstatus_csv_dumper_1096 = new("./chan_status1096.csv");
    fifo_monitor_1096 = new(fifo_csv_dumper_1096,fifo_intf_1096,cstatus_csv_dumper_1096);
    fifo_csv_dumper_1097 = new("./depth1097.csv");
    cstatus_csv_dumper_1097 = new("./chan_status1097.csv");
    fifo_monitor_1097 = new(fifo_csv_dumper_1097,fifo_intf_1097,cstatus_csv_dumper_1097);
    fifo_csv_dumper_1098 = new("./depth1098.csv");
    cstatus_csv_dumper_1098 = new("./chan_status1098.csv");
    fifo_monitor_1098 = new(fifo_csv_dumper_1098,fifo_intf_1098,cstatus_csv_dumper_1098);
    fifo_csv_dumper_1099 = new("./depth1099.csv");
    cstatus_csv_dumper_1099 = new("./chan_status1099.csv");
    fifo_monitor_1099 = new(fifo_csv_dumper_1099,fifo_intf_1099,cstatus_csv_dumper_1099);
    fifo_csv_dumper_1100 = new("./depth1100.csv");
    cstatus_csv_dumper_1100 = new("./chan_status1100.csv");
    fifo_monitor_1100 = new(fifo_csv_dumper_1100,fifo_intf_1100,cstatus_csv_dumper_1100);
    fifo_csv_dumper_1101 = new("./depth1101.csv");
    cstatus_csv_dumper_1101 = new("./chan_status1101.csv");
    fifo_monitor_1101 = new(fifo_csv_dumper_1101,fifo_intf_1101,cstatus_csv_dumper_1101);
    fifo_csv_dumper_1102 = new("./depth1102.csv");
    cstatus_csv_dumper_1102 = new("./chan_status1102.csv");
    fifo_monitor_1102 = new(fifo_csv_dumper_1102,fifo_intf_1102,cstatus_csv_dumper_1102);
    fifo_csv_dumper_1103 = new("./depth1103.csv");
    cstatus_csv_dumper_1103 = new("./chan_status1103.csv");
    fifo_monitor_1103 = new(fifo_csv_dumper_1103,fifo_intf_1103,cstatus_csv_dumper_1103);
    fifo_csv_dumper_1104 = new("./depth1104.csv");
    cstatus_csv_dumper_1104 = new("./chan_status1104.csv");
    fifo_monitor_1104 = new(fifo_csv_dumper_1104,fifo_intf_1104,cstatus_csv_dumper_1104);
    fifo_csv_dumper_1105 = new("./depth1105.csv");
    cstatus_csv_dumper_1105 = new("./chan_status1105.csv");
    fifo_monitor_1105 = new(fifo_csv_dumper_1105,fifo_intf_1105,cstatus_csv_dumper_1105);
    fifo_csv_dumper_1106 = new("./depth1106.csv");
    cstatus_csv_dumper_1106 = new("./chan_status1106.csv");
    fifo_monitor_1106 = new(fifo_csv_dumper_1106,fifo_intf_1106,cstatus_csv_dumper_1106);
    fifo_csv_dumper_1107 = new("./depth1107.csv");
    cstatus_csv_dumper_1107 = new("./chan_status1107.csv");
    fifo_monitor_1107 = new(fifo_csv_dumper_1107,fifo_intf_1107,cstatus_csv_dumper_1107);
    fifo_csv_dumper_1108 = new("./depth1108.csv");
    cstatus_csv_dumper_1108 = new("./chan_status1108.csv");
    fifo_monitor_1108 = new(fifo_csv_dumper_1108,fifo_intf_1108,cstatus_csv_dumper_1108);
    fifo_csv_dumper_1109 = new("./depth1109.csv");
    cstatus_csv_dumper_1109 = new("./chan_status1109.csv");
    fifo_monitor_1109 = new(fifo_csv_dumper_1109,fifo_intf_1109,cstatus_csv_dumper_1109);
    fifo_csv_dumper_1110 = new("./depth1110.csv");
    cstatus_csv_dumper_1110 = new("./chan_status1110.csv");
    fifo_monitor_1110 = new(fifo_csv_dumper_1110,fifo_intf_1110,cstatus_csv_dumper_1110);
    fifo_csv_dumper_1111 = new("./depth1111.csv");
    cstatus_csv_dumper_1111 = new("./chan_status1111.csv");
    fifo_monitor_1111 = new(fifo_csv_dumper_1111,fifo_intf_1111,cstatus_csv_dumper_1111);
    fifo_csv_dumper_1112 = new("./depth1112.csv");
    cstatus_csv_dumper_1112 = new("./chan_status1112.csv");
    fifo_monitor_1112 = new(fifo_csv_dumper_1112,fifo_intf_1112,cstatus_csv_dumper_1112);
    fifo_csv_dumper_1113 = new("./depth1113.csv");
    cstatus_csv_dumper_1113 = new("./chan_status1113.csv");
    fifo_monitor_1113 = new(fifo_csv_dumper_1113,fifo_intf_1113,cstatus_csv_dumper_1113);
    fifo_csv_dumper_1114 = new("./depth1114.csv");
    cstatus_csv_dumper_1114 = new("./chan_status1114.csv");
    fifo_monitor_1114 = new(fifo_csv_dumper_1114,fifo_intf_1114,cstatus_csv_dumper_1114);
    fifo_csv_dumper_1115 = new("./depth1115.csv");
    cstatus_csv_dumper_1115 = new("./chan_status1115.csv");
    fifo_monitor_1115 = new(fifo_csv_dumper_1115,fifo_intf_1115,cstatus_csv_dumper_1115);
    fifo_csv_dumper_1116 = new("./depth1116.csv");
    cstatus_csv_dumper_1116 = new("./chan_status1116.csv");
    fifo_monitor_1116 = new(fifo_csv_dumper_1116,fifo_intf_1116,cstatus_csv_dumper_1116);
    fifo_csv_dumper_1117 = new("./depth1117.csv");
    cstatus_csv_dumper_1117 = new("./chan_status1117.csv");
    fifo_monitor_1117 = new(fifo_csv_dumper_1117,fifo_intf_1117,cstatus_csv_dumper_1117);
    fifo_csv_dumper_1118 = new("./depth1118.csv");
    cstatus_csv_dumper_1118 = new("./chan_status1118.csv");
    fifo_monitor_1118 = new(fifo_csv_dumper_1118,fifo_intf_1118,cstatus_csv_dumper_1118);
    fifo_csv_dumper_1119 = new("./depth1119.csv");
    cstatus_csv_dumper_1119 = new("./chan_status1119.csv");
    fifo_monitor_1119 = new(fifo_csv_dumper_1119,fifo_intf_1119,cstatus_csv_dumper_1119);
    fifo_csv_dumper_1120 = new("./depth1120.csv");
    cstatus_csv_dumper_1120 = new("./chan_status1120.csv");
    fifo_monitor_1120 = new(fifo_csv_dumper_1120,fifo_intf_1120,cstatus_csv_dumper_1120);
    fifo_csv_dumper_1121 = new("./depth1121.csv");
    cstatus_csv_dumper_1121 = new("./chan_status1121.csv");
    fifo_monitor_1121 = new(fifo_csv_dumper_1121,fifo_intf_1121,cstatus_csv_dumper_1121);
    fifo_csv_dumper_1122 = new("./depth1122.csv");
    cstatus_csv_dumper_1122 = new("./chan_status1122.csv");
    fifo_monitor_1122 = new(fifo_csv_dumper_1122,fifo_intf_1122,cstatus_csv_dumper_1122);
    fifo_csv_dumper_1123 = new("./depth1123.csv");
    cstatus_csv_dumper_1123 = new("./chan_status1123.csv");
    fifo_monitor_1123 = new(fifo_csv_dumper_1123,fifo_intf_1123,cstatus_csv_dumper_1123);
    fifo_csv_dumper_1124 = new("./depth1124.csv");
    cstatus_csv_dumper_1124 = new("./chan_status1124.csv");
    fifo_monitor_1124 = new(fifo_csv_dumper_1124,fifo_intf_1124,cstatus_csv_dumper_1124);
    fifo_csv_dumper_1125 = new("./depth1125.csv");
    cstatus_csv_dumper_1125 = new("./chan_status1125.csv");
    fifo_monitor_1125 = new(fifo_csv_dumper_1125,fifo_intf_1125,cstatus_csv_dumper_1125);
    fifo_csv_dumper_1126 = new("./depth1126.csv");
    cstatus_csv_dumper_1126 = new("./chan_status1126.csv");
    fifo_monitor_1126 = new(fifo_csv_dumper_1126,fifo_intf_1126,cstatus_csv_dumper_1126);
    fifo_csv_dumper_1127 = new("./depth1127.csv");
    cstatus_csv_dumper_1127 = new("./chan_status1127.csv");
    fifo_monitor_1127 = new(fifo_csv_dumper_1127,fifo_intf_1127,cstatus_csv_dumper_1127);
    fifo_csv_dumper_1128 = new("./depth1128.csv");
    cstatus_csv_dumper_1128 = new("./chan_status1128.csv");
    fifo_monitor_1128 = new(fifo_csv_dumper_1128,fifo_intf_1128,cstatus_csv_dumper_1128);
    fifo_csv_dumper_1129 = new("./depth1129.csv");
    cstatus_csv_dumper_1129 = new("./chan_status1129.csv");
    fifo_monitor_1129 = new(fifo_csv_dumper_1129,fifo_intf_1129,cstatus_csv_dumper_1129);
    fifo_csv_dumper_1130 = new("./depth1130.csv");
    cstatus_csv_dumper_1130 = new("./chan_status1130.csv");
    fifo_monitor_1130 = new(fifo_csv_dumper_1130,fifo_intf_1130,cstatus_csv_dumper_1130);
    fifo_csv_dumper_1131 = new("./depth1131.csv");
    cstatus_csv_dumper_1131 = new("./chan_status1131.csv");
    fifo_monitor_1131 = new(fifo_csv_dumper_1131,fifo_intf_1131,cstatus_csv_dumper_1131);
    fifo_csv_dumper_1132 = new("./depth1132.csv");
    cstatus_csv_dumper_1132 = new("./chan_status1132.csv");
    fifo_monitor_1132 = new(fifo_csv_dumper_1132,fifo_intf_1132,cstatus_csv_dumper_1132);
    fifo_csv_dumper_1133 = new("./depth1133.csv");
    cstatus_csv_dumper_1133 = new("./chan_status1133.csv");
    fifo_monitor_1133 = new(fifo_csv_dumper_1133,fifo_intf_1133,cstatus_csv_dumper_1133);
    fifo_csv_dumper_1134 = new("./depth1134.csv");
    cstatus_csv_dumper_1134 = new("./chan_status1134.csv");
    fifo_monitor_1134 = new(fifo_csv_dumper_1134,fifo_intf_1134,cstatus_csv_dumper_1134);
    fifo_csv_dumper_1135 = new("./depth1135.csv");
    cstatus_csv_dumper_1135 = new("./chan_status1135.csv");
    fifo_monitor_1135 = new(fifo_csv_dumper_1135,fifo_intf_1135,cstatus_csv_dumper_1135);
    fifo_csv_dumper_1136 = new("./depth1136.csv");
    cstatus_csv_dumper_1136 = new("./chan_status1136.csv");
    fifo_monitor_1136 = new(fifo_csv_dumper_1136,fifo_intf_1136,cstatus_csv_dumper_1136);
    fifo_csv_dumper_1137 = new("./depth1137.csv");
    cstatus_csv_dumper_1137 = new("./chan_status1137.csv");
    fifo_monitor_1137 = new(fifo_csv_dumper_1137,fifo_intf_1137,cstatus_csv_dumper_1137);
    fifo_csv_dumper_1138 = new("./depth1138.csv");
    cstatus_csv_dumper_1138 = new("./chan_status1138.csv");
    fifo_monitor_1138 = new(fifo_csv_dumper_1138,fifo_intf_1138,cstatus_csv_dumper_1138);
    fifo_csv_dumper_1139 = new("./depth1139.csv");
    cstatus_csv_dumper_1139 = new("./chan_status1139.csv");
    fifo_monitor_1139 = new(fifo_csv_dumper_1139,fifo_intf_1139,cstatus_csv_dumper_1139);
    fifo_csv_dumper_1140 = new("./depth1140.csv");
    cstatus_csv_dumper_1140 = new("./chan_status1140.csv");
    fifo_monitor_1140 = new(fifo_csv_dumper_1140,fifo_intf_1140,cstatus_csv_dumper_1140);
    fifo_csv_dumper_1141 = new("./depth1141.csv");
    cstatus_csv_dumper_1141 = new("./chan_status1141.csv");
    fifo_monitor_1141 = new(fifo_csv_dumper_1141,fifo_intf_1141,cstatus_csv_dumper_1141);
    fifo_csv_dumper_1142 = new("./depth1142.csv");
    cstatus_csv_dumper_1142 = new("./chan_status1142.csv");
    fifo_monitor_1142 = new(fifo_csv_dumper_1142,fifo_intf_1142,cstatus_csv_dumper_1142);
    fifo_csv_dumper_1143 = new("./depth1143.csv");
    cstatus_csv_dumper_1143 = new("./chan_status1143.csv");
    fifo_monitor_1143 = new(fifo_csv_dumper_1143,fifo_intf_1143,cstatus_csv_dumper_1143);
    fifo_csv_dumper_1144 = new("./depth1144.csv");
    cstatus_csv_dumper_1144 = new("./chan_status1144.csv");
    fifo_monitor_1144 = new(fifo_csv_dumper_1144,fifo_intf_1144,cstatus_csv_dumper_1144);
    fifo_csv_dumper_1145 = new("./depth1145.csv");
    cstatus_csv_dumper_1145 = new("./chan_status1145.csv");
    fifo_monitor_1145 = new(fifo_csv_dumper_1145,fifo_intf_1145,cstatus_csv_dumper_1145);
    fifo_csv_dumper_1146 = new("./depth1146.csv");
    cstatus_csv_dumper_1146 = new("./chan_status1146.csv");
    fifo_monitor_1146 = new(fifo_csv_dumper_1146,fifo_intf_1146,cstatus_csv_dumper_1146);
    fifo_csv_dumper_1147 = new("./depth1147.csv");
    cstatus_csv_dumper_1147 = new("./chan_status1147.csv");
    fifo_monitor_1147 = new(fifo_csv_dumper_1147,fifo_intf_1147,cstatus_csv_dumper_1147);
    fifo_csv_dumper_1148 = new("./depth1148.csv");
    cstatus_csv_dumper_1148 = new("./chan_status1148.csv");
    fifo_monitor_1148 = new(fifo_csv_dumper_1148,fifo_intf_1148,cstatus_csv_dumper_1148);
    fifo_csv_dumper_1149 = new("./depth1149.csv");
    cstatus_csv_dumper_1149 = new("./chan_status1149.csv");
    fifo_monitor_1149 = new(fifo_csv_dumper_1149,fifo_intf_1149,cstatus_csv_dumper_1149);
    fifo_csv_dumper_1150 = new("./depth1150.csv");
    cstatus_csv_dumper_1150 = new("./chan_status1150.csv");
    fifo_monitor_1150 = new(fifo_csv_dumper_1150,fifo_intf_1150,cstatus_csv_dumper_1150);
    fifo_csv_dumper_1151 = new("./depth1151.csv");
    cstatus_csv_dumper_1151 = new("./chan_status1151.csv");
    fifo_monitor_1151 = new(fifo_csv_dumper_1151,fifo_intf_1151,cstatus_csv_dumper_1151);
    fifo_csv_dumper_1152 = new("./depth1152.csv");
    cstatus_csv_dumper_1152 = new("./chan_status1152.csv");
    fifo_monitor_1152 = new(fifo_csv_dumper_1152,fifo_intf_1152,cstatus_csv_dumper_1152);
    fifo_csv_dumper_1153 = new("./depth1153.csv");
    cstatus_csv_dumper_1153 = new("./chan_status1153.csv");
    fifo_monitor_1153 = new(fifo_csv_dumper_1153,fifo_intf_1153,cstatus_csv_dumper_1153);
    fifo_csv_dumper_1154 = new("./depth1154.csv");
    cstatus_csv_dumper_1154 = new("./chan_status1154.csv");
    fifo_monitor_1154 = new(fifo_csv_dumper_1154,fifo_intf_1154,cstatus_csv_dumper_1154);
    fifo_csv_dumper_1155 = new("./depth1155.csv");
    cstatus_csv_dumper_1155 = new("./chan_status1155.csv");
    fifo_monitor_1155 = new(fifo_csv_dumper_1155,fifo_intf_1155,cstatus_csv_dumper_1155);
    fifo_csv_dumper_1156 = new("./depth1156.csv");
    cstatus_csv_dumper_1156 = new("./chan_status1156.csv");
    fifo_monitor_1156 = new(fifo_csv_dumper_1156,fifo_intf_1156,cstatus_csv_dumper_1156);
    fifo_csv_dumper_1157 = new("./depth1157.csv");
    cstatus_csv_dumper_1157 = new("./chan_status1157.csv");
    fifo_monitor_1157 = new(fifo_csv_dumper_1157,fifo_intf_1157,cstatus_csv_dumper_1157);
    fifo_csv_dumper_1158 = new("./depth1158.csv");
    cstatus_csv_dumper_1158 = new("./chan_status1158.csv");
    fifo_monitor_1158 = new(fifo_csv_dumper_1158,fifo_intf_1158,cstatus_csv_dumper_1158);
    fifo_csv_dumper_1159 = new("./depth1159.csv");
    cstatus_csv_dumper_1159 = new("./chan_status1159.csv");
    fifo_monitor_1159 = new(fifo_csv_dumper_1159,fifo_intf_1159,cstatus_csv_dumper_1159);
    fifo_csv_dumper_1160 = new("./depth1160.csv");
    cstatus_csv_dumper_1160 = new("./chan_status1160.csv");
    fifo_monitor_1160 = new(fifo_csv_dumper_1160,fifo_intf_1160,cstatus_csv_dumper_1160);
    fifo_csv_dumper_1161 = new("./depth1161.csv");
    cstatus_csv_dumper_1161 = new("./chan_status1161.csv");
    fifo_monitor_1161 = new(fifo_csv_dumper_1161,fifo_intf_1161,cstatus_csv_dumper_1161);
    fifo_csv_dumper_1162 = new("./depth1162.csv");
    cstatus_csv_dumper_1162 = new("./chan_status1162.csv");
    fifo_monitor_1162 = new(fifo_csv_dumper_1162,fifo_intf_1162,cstatus_csv_dumper_1162);
    fifo_csv_dumper_1163 = new("./depth1163.csv");
    cstatus_csv_dumper_1163 = new("./chan_status1163.csv");
    fifo_monitor_1163 = new(fifo_csv_dumper_1163,fifo_intf_1163,cstatus_csv_dumper_1163);
    fifo_csv_dumper_1164 = new("./depth1164.csv");
    cstatus_csv_dumper_1164 = new("./chan_status1164.csv");
    fifo_monitor_1164 = new(fifo_csv_dumper_1164,fifo_intf_1164,cstatus_csv_dumper_1164);
    fifo_csv_dumper_1165 = new("./depth1165.csv");
    cstatus_csv_dumper_1165 = new("./chan_status1165.csv");
    fifo_monitor_1165 = new(fifo_csv_dumper_1165,fifo_intf_1165,cstatus_csv_dumper_1165);
    fifo_csv_dumper_1166 = new("./depth1166.csv");
    cstatus_csv_dumper_1166 = new("./chan_status1166.csv");
    fifo_monitor_1166 = new(fifo_csv_dumper_1166,fifo_intf_1166,cstatus_csv_dumper_1166);
    fifo_csv_dumper_1167 = new("./depth1167.csv");
    cstatus_csv_dumper_1167 = new("./chan_status1167.csv");
    fifo_monitor_1167 = new(fifo_csv_dumper_1167,fifo_intf_1167,cstatus_csv_dumper_1167);
    fifo_csv_dumper_1168 = new("./depth1168.csv");
    cstatus_csv_dumper_1168 = new("./chan_status1168.csv");
    fifo_monitor_1168 = new(fifo_csv_dumper_1168,fifo_intf_1168,cstatus_csv_dumper_1168);
    fifo_csv_dumper_1169 = new("./depth1169.csv");
    cstatus_csv_dumper_1169 = new("./chan_status1169.csv");
    fifo_monitor_1169 = new(fifo_csv_dumper_1169,fifo_intf_1169,cstatus_csv_dumper_1169);
    fifo_csv_dumper_1170 = new("./depth1170.csv");
    cstatus_csv_dumper_1170 = new("./chan_status1170.csv");
    fifo_monitor_1170 = new(fifo_csv_dumper_1170,fifo_intf_1170,cstatus_csv_dumper_1170);
    fifo_csv_dumper_1171 = new("./depth1171.csv");
    cstatus_csv_dumper_1171 = new("./chan_status1171.csv");
    fifo_monitor_1171 = new(fifo_csv_dumper_1171,fifo_intf_1171,cstatus_csv_dumper_1171);
    fifo_csv_dumper_1172 = new("./depth1172.csv");
    cstatus_csv_dumper_1172 = new("./chan_status1172.csv");
    fifo_monitor_1172 = new(fifo_csv_dumper_1172,fifo_intf_1172,cstatus_csv_dumper_1172);
    fifo_csv_dumper_1173 = new("./depth1173.csv");
    cstatus_csv_dumper_1173 = new("./chan_status1173.csv");
    fifo_monitor_1173 = new(fifo_csv_dumper_1173,fifo_intf_1173,cstatus_csv_dumper_1173);
    fifo_csv_dumper_1174 = new("./depth1174.csv");
    cstatus_csv_dumper_1174 = new("./chan_status1174.csv");
    fifo_monitor_1174 = new(fifo_csv_dumper_1174,fifo_intf_1174,cstatus_csv_dumper_1174);
    fifo_csv_dumper_1175 = new("./depth1175.csv");
    cstatus_csv_dumper_1175 = new("./chan_status1175.csv");
    fifo_monitor_1175 = new(fifo_csv_dumper_1175,fifo_intf_1175,cstatus_csv_dumper_1175);
    fifo_csv_dumper_1176 = new("./depth1176.csv");
    cstatus_csv_dumper_1176 = new("./chan_status1176.csv");
    fifo_monitor_1176 = new(fifo_csv_dumper_1176,fifo_intf_1176,cstatus_csv_dumper_1176);
    fifo_csv_dumper_1177 = new("./depth1177.csv");
    cstatus_csv_dumper_1177 = new("./chan_status1177.csv");
    fifo_monitor_1177 = new(fifo_csv_dumper_1177,fifo_intf_1177,cstatus_csv_dumper_1177);
    fifo_csv_dumper_1178 = new("./depth1178.csv");
    cstatus_csv_dumper_1178 = new("./chan_status1178.csv");
    fifo_monitor_1178 = new(fifo_csv_dumper_1178,fifo_intf_1178,cstatus_csv_dumper_1178);
    fifo_csv_dumper_1179 = new("./depth1179.csv");
    cstatus_csv_dumper_1179 = new("./chan_status1179.csv");
    fifo_monitor_1179 = new(fifo_csv_dumper_1179,fifo_intf_1179,cstatus_csv_dumper_1179);
    fifo_csv_dumper_1180 = new("./depth1180.csv");
    cstatus_csv_dumper_1180 = new("./chan_status1180.csv");
    fifo_monitor_1180 = new(fifo_csv_dumper_1180,fifo_intf_1180,cstatus_csv_dumper_1180);
    fifo_csv_dumper_1181 = new("./depth1181.csv");
    cstatus_csv_dumper_1181 = new("./chan_status1181.csv");
    fifo_monitor_1181 = new(fifo_csv_dumper_1181,fifo_intf_1181,cstatus_csv_dumper_1181);
    fifo_csv_dumper_1182 = new("./depth1182.csv");
    cstatus_csv_dumper_1182 = new("./chan_status1182.csv");
    fifo_monitor_1182 = new(fifo_csv_dumper_1182,fifo_intf_1182,cstatus_csv_dumper_1182);
    fifo_csv_dumper_1183 = new("./depth1183.csv");
    cstatus_csv_dumper_1183 = new("./chan_status1183.csv");
    fifo_monitor_1183 = new(fifo_csv_dumper_1183,fifo_intf_1183,cstatus_csv_dumper_1183);
    fifo_csv_dumper_1184 = new("./depth1184.csv");
    cstatus_csv_dumper_1184 = new("./chan_status1184.csv");
    fifo_monitor_1184 = new(fifo_csv_dumper_1184,fifo_intf_1184,cstatus_csv_dumper_1184);
    fifo_csv_dumper_1185 = new("./depth1185.csv");
    cstatus_csv_dumper_1185 = new("./chan_status1185.csv");
    fifo_monitor_1185 = new(fifo_csv_dumper_1185,fifo_intf_1185,cstatus_csv_dumper_1185);
    fifo_csv_dumper_1186 = new("./depth1186.csv");
    cstatus_csv_dumper_1186 = new("./chan_status1186.csv");
    fifo_monitor_1186 = new(fifo_csv_dumper_1186,fifo_intf_1186,cstatus_csv_dumper_1186);
    fifo_csv_dumper_1187 = new("./depth1187.csv");
    cstatus_csv_dumper_1187 = new("./chan_status1187.csv");
    fifo_monitor_1187 = new(fifo_csv_dumper_1187,fifo_intf_1187,cstatus_csv_dumper_1187);
    fifo_csv_dumper_1188 = new("./depth1188.csv");
    cstatus_csv_dumper_1188 = new("./chan_status1188.csv");
    fifo_monitor_1188 = new(fifo_csv_dumper_1188,fifo_intf_1188,cstatus_csv_dumper_1188);
    fifo_csv_dumper_1189 = new("./depth1189.csv");
    cstatus_csv_dumper_1189 = new("./chan_status1189.csv");
    fifo_monitor_1189 = new(fifo_csv_dumper_1189,fifo_intf_1189,cstatus_csv_dumper_1189);
    fifo_csv_dumper_1190 = new("./depth1190.csv");
    cstatus_csv_dumper_1190 = new("./chan_status1190.csv");
    fifo_monitor_1190 = new(fifo_csv_dumper_1190,fifo_intf_1190,cstatus_csv_dumper_1190);
    fifo_csv_dumper_1191 = new("./depth1191.csv");
    cstatus_csv_dumper_1191 = new("./chan_status1191.csv");
    fifo_monitor_1191 = new(fifo_csv_dumper_1191,fifo_intf_1191,cstatus_csv_dumper_1191);
    fifo_csv_dumper_1192 = new("./depth1192.csv");
    cstatus_csv_dumper_1192 = new("./chan_status1192.csv");
    fifo_monitor_1192 = new(fifo_csv_dumper_1192,fifo_intf_1192,cstatus_csv_dumper_1192);
    fifo_csv_dumper_1193 = new("./depth1193.csv");
    cstatus_csv_dumper_1193 = new("./chan_status1193.csv");
    fifo_monitor_1193 = new(fifo_csv_dumper_1193,fifo_intf_1193,cstatus_csv_dumper_1193);
    fifo_csv_dumper_1194 = new("./depth1194.csv");
    cstatus_csv_dumper_1194 = new("./chan_status1194.csv");
    fifo_monitor_1194 = new(fifo_csv_dumper_1194,fifo_intf_1194,cstatus_csv_dumper_1194);
    fifo_csv_dumper_1195 = new("./depth1195.csv");
    cstatus_csv_dumper_1195 = new("./chan_status1195.csv");
    fifo_monitor_1195 = new(fifo_csv_dumper_1195,fifo_intf_1195,cstatus_csv_dumper_1195);
    fifo_csv_dumper_1196 = new("./depth1196.csv");
    cstatus_csv_dumper_1196 = new("./chan_status1196.csv");
    fifo_monitor_1196 = new(fifo_csv_dumper_1196,fifo_intf_1196,cstatus_csv_dumper_1196);
    fifo_csv_dumper_1197 = new("./depth1197.csv");
    cstatus_csv_dumper_1197 = new("./chan_status1197.csv");
    fifo_monitor_1197 = new(fifo_csv_dumper_1197,fifo_intf_1197,cstatus_csv_dumper_1197);
    fifo_csv_dumper_1198 = new("./depth1198.csv");
    cstatus_csv_dumper_1198 = new("./chan_status1198.csv");
    fifo_monitor_1198 = new(fifo_csv_dumper_1198,fifo_intf_1198,cstatus_csv_dumper_1198);
    fifo_csv_dumper_1199 = new("./depth1199.csv");
    cstatus_csv_dumper_1199 = new("./chan_status1199.csv");
    fifo_monitor_1199 = new(fifo_csv_dumper_1199,fifo_intf_1199,cstatus_csv_dumper_1199);
    fifo_csv_dumper_1200 = new("./depth1200.csv");
    cstatus_csv_dumper_1200 = new("./chan_status1200.csv");
    fifo_monitor_1200 = new(fifo_csv_dumper_1200,fifo_intf_1200,cstatus_csv_dumper_1200);
    fifo_csv_dumper_1201 = new("./depth1201.csv");
    cstatus_csv_dumper_1201 = new("./chan_status1201.csv");
    fifo_monitor_1201 = new(fifo_csv_dumper_1201,fifo_intf_1201,cstatus_csv_dumper_1201);
    fifo_csv_dumper_1202 = new("./depth1202.csv");
    cstatus_csv_dumper_1202 = new("./chan_status1202.csv");
    fifo_monitor_1202 = new(fifo_csv_dumper_1202,fifo_intf_1202,cstatus_csv_dumper_1202);
    fifo_csv_dumper_1203 = new("./depth1203.csv");
    cstatus_csv_dumper_1203 = new("./chan_status1203.csv");
    fifo_monitor_1203 = new(fifo_csv_dumper_1203,fifo_intf_1203,cstatus_csv_dumper_1203);
    fifo_csv_dumper_1204 = new("./depth1204.csv");
    cstatus_csv_dumper_1204 = new("./chan_status1204.csv");
    fifo_monitor_1204 = new(fifo_csv_dumper_1204,fifo_intf_1204,cstatus_csv_dumper_1204);
    fifo_csv_dumper_1205 = new("./depth1205.csv");
    cstatus_csv_dumper_1205 = new("./chan_status1205.csv");
    fifo_monitor_1205 = new(fifo_csv_dumper_1205,fifo_intf_1205,cstatus_csv_dumper_1205);
    fifo_csv_dumper_1206 = new("./depth1206.csv");
    cstatus_csv_dumper_1206 = new("./chan_status1206.csv");
    fifo_monitor_1206 = new(fifo_csv_dumper_1206,fifo_intf_1206,cstatus_csv_dumper_1206);
    fifo_csv_dumper_1207 = new("./depth1207.csv");
    cstatus_csv_dumper_1207 = new("./chan_status1207.csv");
    fifo_monitor_1207 = new(fifo_csv_dumper_1207,fifo_intf_1207,cstatus_csv_dumper_1207);
    fifo_csv_dumper_1208 = new("./depth1208.csv");
    cstatus_csv_dumper_1208 = new("./chan_status1208.csv");
    fifo_monitor_1208 = new(fifo_csv_dumper_1208,fifo_intf_1208,cstatus_csv_dumper_1208);
    fifo_csv_dumper_1209 = new("./depth1209.csv");
    cstatus_csv_dumper_1209 = new("./chan_status1209.csv");
    fifo_monitor_1209 = new(fifo_csv_dumper_1209,fifo_intf_1209,cstatus_csv_dumper_1209);
    fifo_csv_dumper_1210 = new("./depth1210.csv");
    cstatus_csv_dumper_1210 = new("./chan_status1210.csv");
    fifo_monitor_1210 = new(fifo_csv_dumper_1210,fifo_intf_1210,cstatus_csv_dumper_1210);
    fifo_csv_dumper_1211 = new("./depth1211.csv");
    cstatus_csv_dumper_1211 = new("./chan_status1211.csv");
    fifo_monitor_1211 = new(fifo_csv_dumper_1211,fifo_intf_1211,cstatus_csv_dumper_1211);
    fifo_csv_dumper_1212 = new("./depth1212.csv");
    cstatus_csv_dumper_1212 = new("./chan_status1212.csv");
    fifo_monitor_1212 = new(fifo_csv_dumper_1212,fifo_intf_1212,cstatus_csv_dumper_1212);
    fifo_csv_dumper_1213 = new("./depth1213.csv");
    cstatus_csv_dumper_1213 = new("./chan_status1213.csv");
    fifo_monitor_1213 = new(fifo_csv_dumper_1213,fifo_intf_1213,cstatus_csv_dumper_1213);
    fifo_csv_dumper_1214 = new("./depth1214.csv");
    cstatus_csv_dumper_1214 = new("./chan_status1214.csv");
    fifo_monitor_1214 = new(fifo_csv_dumper_1214,fifo_intf_1214,cstatus_csv_dumper_1214);
    fifo_csv_dumper_1215 = new("./depth1215.csv");
    cstatus_csv_dumper_1215 = new("./chan_status1215.csv");
    fifo_monitor_1215 = new(fifo_csv_dumper_1215,fifo_intf_1215,cstatus_csv_dumper_1215);
    fifo_csv_dumper_1216 = new("./depth1216.csv");
    cstatus_csv_dumper_1216 = new("./chan_status1216.csv");
    fifo_monitor_1216 = new(fifo_csv_dumper_1216,fifo_intf_1216,cstatus_csv_dumper_1216);
    fifo_csv_dumper_1217 = new("./depth1217.csv");
    cstatus_csv_dumper_1217 = new("./chan_status1217.csv");
    fifo_monitor_1217 = new(fifo_csv_dumper_1217,fifo_intf_1217,cstatus_csv_dumper_1217);
    fifo_csv_dumper_1218 = new("./depth1218.csv");
    cstatus_csv_dumper_1218 = new("./chan_status1218.csv");
    fifo_monitor_1218 = new(fifo_csv_dumper_1218,fifo_intf_1218,cstatus_csv_dumper_1218);
    fifo_csv_dumper_1219 = new("./depth1219.csv");
    cstatus_csv_dumper_1219 = new("./chan_status1219.csv");
    fifo_monitor_1219 = new(fifo_csv_dumper_1219,fifo_intf_1219,cstatus_csv_dumper_1219);
    fifo_csv_dumper_1220 = new("./depth1220.csv");
    cstatus_csv_dumper_1220 = new("./chan_status1220.csv");
    fifo_monitor_1220 = new(fifo_csv_dumper_1220,fifo_intf_1220,cstatus_csv_dumper_1220);
    fifo_csv_dumper_1221 = new("./depth1221.csv");
    cstatus_csv_dumper_1221 = new("./chan_status1221.csv");
    fifo_monitor_1221 = new(fifo_csv_dumper_1221,fifo_intf_1221,cstatus_csv_dumper_1221);
    fifo_csv_dumper_1222 = new("./depth1222.csv");
    cstatus_csv_dumper_1222 = new("./chan_status1222.csv");
    fifo_monitor_1222 = new(fifo_csv_dumper_1222,fifo_intf_1222,cstatus_csv_dumper_1222);
    fifo_csv_dumper_1223 = new("./depth1223.csv");
    cstatus_csv_dumper_1223 = new("./chan_status1223.csv");
    fifo_monitor_1223 = new(fifo_csv_dumper_1223,fifo_intf_1223,cstatus_csv_dumper_1223);
    fifo_csv_dumper_1224 = new("./depth1224.csv");
    cstatus_csv_dumper_1224 = new("./chan_status1224.csv");
    fifo_monitor_1224 = new(fifo_csv_dumper_1224,fifo_intf_1224,cstatus_csv_dumper_1224);
    fifo_csv_dumper_1225 = new("./depth1225.csv");
    cstatus_csv_dumper_1225 = new("./chan_status1225.csv");
    fifo_monitor_1225 = new(fifo_csv_dumper_1225,fifo_intf_1225,cstatus_csv_dumper_1225);
    fifo_csv_dumper_1226 = new("./depth1226.csv");
    cstatus_csv_dumper_1226 = new("./chan_status1226.csv");
    fifo_monitor_1226 = new(fifo_csv_dumper_1226,fifo_intf_1226,cstatus_csv_dumper_1226);
    fifo_csv_dumper_1227 = new("./depth1227.csv");
    cstatus_csv_dumper_1227 = new("./chan_status1227.csv");
    fifo_monitor_1227 = new(fifo_csv_dumper_1227,fifo_intf_1227,cstatus_csv_dumper_1227);
    fifo_csv_dumper_1228 = new("./depth1228.csv");
    cstatus_csv_dumper_1228 = new("./chan_status1228.csv");
    fifo_monitor_1228 = new(fifo_csv_dumper_1228,fifo_intf_1228,cstatus_csv_dumper_1228);
    fifo_csv_dumper_1229 = new("./depth1229.csv");
    cstatus_csv_dumper_1229 = new("./chan_status1229.csv");
    fifo_monitor_1229 = new(fifo_csv_dumper_1229,fifo_intf_1229,cstatus_csv_dumper_1229);
    fifo_csv_dumper_1230 = new("./depth1230.csv");
    cstatus_csv_dumper_1230 = new("./chan_status1230.csv");
    fifo_monitor_1230 = new(fifo_csv_dumper_1230,fifo_intf_1230,cstatus_csv_dumper_1230);
    fifo_csv_dumper_1231 = new("./depth1231.csv");
    cstatus_csv_dumper_1231 = new("./chan_status1231.csv");
    fifo_monitor_1231 = new(fifo_csv_dumper_1231,fifo_intf_1231,cstatus_csv_dumper_1231);
    fifo_csv_dumper_1232 = new("./depth1232.csv");
    cstatus_csv_dumper_1232 = new("./chan_status1232.csv");
    fifo_monitor_1232 = new(fifo_csv_dumper_1232,fifo_intf_1232,cstatus_csv_dumper_1232);
    fifo_csv_dumper_1233 = new("./depth1233.csv");
    cstatus_csv_dumper_1233 = new("./chan_status1233.csv");
    fifo_monitor_1233 = new(fifo_csv_dumper_1233,fifo_intf_1233,cstatus_csv_dumper_1233);
    fifo_csv_dumper_1234 = new("./depth1234.csv");
    cstatus_csv_dumper_1234 = new("./chan_status1234.csv");
    fifo_monitor_1234 = new(fifo_csv_dumper_1234,fifo_intf_1234,cstatus_csv_dumper_1234);
    fifo_csv_dumper_1235 = new("./depth1235.csv");
    cstatus_csv_dumper_1235 = new("./chan_status1235.csv");
    fifo_monitor_1235 = new(fifo_csv_dumper_1235,fifo_intf_1235,cstatus_csv_dumper_1235);
    fifo_csv_dumper_1236 = new("./depth1236.csv");
    cstatus_csv_dumper_1236 = new("./chan_status1236.csv");
    fifo_monitor_1236 = new(fifo_csv_dumper_1236,fifo_intf_1236,cstatus_csv_dumper_1236);
    fifo_csv_dumper_1237 = new("./depth1237.csv");
    cstatus_csv_dumper_1237 = new("./chan_status1237.csv");
    fifo_monitor_1237 = new(fifo_csv_dumper_1237,fifo_intf_1237,cstatus_csv_dumper_1237);
    fifo_csv_dumper_1238 = new("./depth1238.csv");
    cstatus_csv_dumper_1238 = new("./chan_status1238.csv");
    fifo_monitor_1238 = new(fifo_csv_dumper_1238,fifo_intf_1238,cstatus_csv_dumper_1238);
    fifo_csv_dumper_1239 = new("./depth1239.csv");
    cstatus_csv_dumper_1239 = new("./chan_status1239.csv");
    fifo_monitor_1239 = new(fifo_csv_dumper_1239,fifo_intf_1239,cstatus_csv_dumper_1239);
    fifo_csv_dumper_1240 = new("./depth1240.csv");
    cstatus_csv_dumper_1240 = new("./chan_status1240.csv");
    fifo_monitor_1240 = new(fifo_csv_dumper_1240,fifo_intf_1240,cstatus_csv_dumper_1240);
    fifo_csv_dumper_1241 = new("./depth1241.csv");
    cstatus_csv_dumper_1241 = new("./chan_status1241.csv");
    fifo_monitor_1241 = new(fifo_csv_dumper_1241,fifo_intf_1241,cstatus_csv_dumper_1241);
    fifo_csv_dumper_1242 = new("./depth1242.csv");
    cstatus_csv_dumper_1242 = new("./chan_status1242.csv");
    fifo_monitor_1242 = new(fifo_csv_dumper_1242,fifo_intf_1242,cstatus_csv_dumper_1242);
    fifo_csv_dumper_1243 = new("./depth1243.csv");
    cstatus_csv_dumper_1243 = new("./chan_status1243.csv");
    fifo_monitor_1243 = new(fifo_csv_dumper_1243,fifo_intf_1243,cstatus_csv_dumper_1243);
    fifo_csv_dumper_1244 = new("./depth1244.csv");
    cstatus_csv_dumper_1244 = new("./chan_status1244.csv");
    fifo_monitor_1244 = new(fifo_csv_dumper_1244,fifo_intf_1244,cstatus_csv_dumper_1244);
    fifo_csv_dumper_1245 = new("./depth1245.csv");
    cstatus_csv_dumper_1245 = new("./chan_status1245.csv");
    fifo_monitor_1245 = new(fifo_csv_dumper_1245,fifo_intf_1245,cstatus_csv_dumper_1245);
    fifo_csv_dumper_1246 = new("./depth1246.csv");
    cstatus_csv_dumper_1246 = new("./chan_status1246.csv");
    fifo_monitor_1246 = new(fifo_csv_dumper_1246,fifo_intf_1246,cstatus_csv_dumper_1246);
    fifo_csv_dumper_1247 = new("./depth1247.csv");
    cstatus_csv_dumper_1247 = new("./chan_status1247.csv");
    fifo_monitor_1247 = new(fifo_csv_dumper_1247,fifo_intf_1247,cstatus_csv_dumper_1247);
    fifo_csv_dumper_1248 = new("./depth1248.csv");
    cstatus_csv_dumper_1248 = new("./chan_status1248.csv");
    fifo_monitor_1248 = new(fifo_csv_dumper_1248,fifo_intf_1248,cstatus_csv_dumper_1248);
    fifo_csv_dumper_1249 = new("./depth1249.csv");
    cstatus_csv_dumper_1249 = new("./chan_status1249.csv");
    fifo_monitor_1249 = new(fifo_csv_dumper_1249,fifo_intf_1249,cstatus_csv_dumper_1249);
    fifo_csv_dumper_1250 = new("./depth1250.csv");
    cstatus_csv_dumper_1250 = new("./chan_status1250.csv");
    fifo_monitor_1250 = new(fifo_csv_dumper_1250,fifo_intf_1250,cstatus_csv_dumper_1250);
    fifo_csv_dumper_1251 = new("./depth1251.csv");
    cstatus_csv_dumper_1251 = new("./chan_status1251.csv");
    fifo_monitor_1251 = new(fifo_csv_dumper_1251,fifo_intf_1251,cstatus_csv_dumper_1251);
    fifo_csv_dumper_1252 = new("./depth1252.csv");
    cstatus_csv_dumper_1252 = new("./chan_status1252.csv");
    fifo_monitor_1252 = new(fifo_csv_dumper_1252,fifo_intf_1252,cstatus_csv_dumper_1252);
    fifo_csv_dumper_1253 = new("./depth1253.csv");
    cstatus_csv_dumper_1253 = new("./chan_status1253.csv");
    fifo_monitor_1253 = new(fifo_csv_dumper_1253,fifo_intf_1253,cstatus_csv_dumper_1253);
    fifo_csv_dumper_1254 = new("./depth1254.csv");
    cstatus_csv_dumper_1254 = new("./chan_status1254.csv");
    fifo_monitor_1254 = new(fifo_csv_dumper_1254,fifo_intf_1254,cstatus_csv_dumper_1254);
    fifo_csv_dumper_1255 = new("./depth1255.csv");
    cstatus_csv_dumper_1255 = new("./chan_status1255.csv");
    fifo_monitor_1255 = new(fifo_csv_dumper_1255,fifo_intf_1255,cstatus_csv_dumper_1255);
    fifo_csv_dumper_1256 = new("./depth1256.csv");
    cstatus_csv_dumper_1256 = new("./chan_status1256.csv");
    fifo_monitor_1256 = new(fifo_csv_dumper_1256,fifo_intf_1256,cstatus_csv_dumper_1256);
    fifo_csv_dumper_1257 = new("./depth1257.csv");
    cstatus_csv_dumper_1257 = new("./chan_status1257.csv");
    fifo_monitor_1257 = new(fifo_csv_dumper_1257,fifo_intf_1257,cstatus_csv_dumper_1257);
    fifo_csv_dumper_1258 = new("./depth1258.csv");
    cstatus_csv_dumper_1258 = new("./chan_status1258.csv");
    fifo_monitor_1258 = new(fifo_csv_dumper_1258,fifo_intf_1258,cstatus_csv_dumper_1258);
    fifo_csv_dumper_1259 = new("./depth1259.csv");
    cstatus_csv_dumper_1259 = new("./chan_status1259.csv");
    fifo_monitor_1259 = new(fifo_csv_dumper_1259,fifo_intf_1259,cstatus_csv_dumper_1259);
    fifo_csv_dumper_1260 = new("./depth1260.csv");
    cstatus_csv_dumper_1260 = new("./chan_status1260.csv");
    fifo_monitor_1260 = new(fifo_csv_dumper_1260,fifo_intf_1260,cstatus_csv_dumper_1260);
    fifo_csv_dumper_1261 = new("./depth1261.csv");
    cstatus_csv_dumper_1261 = new("./chan_status1261.csv");
    fifo_monitor_1261 = new(fifo_csv_dumper_1261,fifo_intf_1261,cstatus_csv_dumper_1261);
    fifo_csv_dumper_1262 = new("./depth1262.csv");
    cstatus_csv_dumper_1262 = new("./chan_status1262.csv");
    fifo_monitor_1262 = new(fifo_csv_dumper_1262,fifo_intf_1262,cstatus_csv_dumper_1262);
    fifo_csv_dumper_1263 = new("./depth1263.csv");
    cstatus_csv_dumper_1263 = new("./chan_status1263.csv");
    fifo_monitor_1263 = new(fifo_csv_dumper_1263,fifo_intf_1263,cstatus_csv_dumper_1263);
    fifo_csv_dumper_1264 = new("./depth1264.csv");
    cstatus_csv_dumper_1264 = new("./chan_status1264.csv");
    fifo_monitor_1264 = new(fifo_csv_dumper_1264,fifo_intf_1264,cstatus_csv_dumper_1264);
    fifo_csv_dumper_1265 = new("./depth1265.csv");
    cstatus_csv_dumper_1265 = new("./chan_status1265.csv");
    fifo_monitor_1265 = new(fifo_csv_dumper_1265,fifo_intf_1265,cstatus_csv_dumper_1265);
    fifo_csv_dumper_1266 = new("./depth1266.csv");
    cstatus_csv_dumper_1266 = new("./chan_status1266.csv");
    fifo_monitor_1266 = new(fifo_csv_dumper_1266,fifo_intf_1266,cstatus_csv_dumper_1266);
    fifo_csv_dumper_1267 = new("./depth1267.csv");
    cstatus_csv_dumper_1267 = new("./chan_status1267.csv");
    fifo_monitor_1267 = new(fifo_csv_dumper_1267,fifo_intf_1267,cstatus_csv_dumper_1267);
    fifo_csv_dumper_1268 = new("./depth1268.csv");
    cstatus_csv_dumper_1268 = new("./chan_status1268.csv");
    fifo_monitor_1268 = new(fifo_csv_dumper_1268,fifo_intf_1268,cstatus_csv_dumper_1268);
    fifo_csv_dumper_1269 = new("./depth1269.csv");
    cstatus_csv_dumper_1269 = new("./chan_status1269.csv");
    fifo_monitor_1269 = new(fifo_csv_dumper_1269,fifo_intf_1269,cstatus_csv_dumper_1269);
    fifo_csv_dumper_1270 = new("./depth1270.csv");
    cstatus_csv_dumper_1270 = new("./chan_status1270.csv");
    fifo_monitor_1270 = new(fifo_csv_dumper_1270,fifo_intf_1270,cstatus_csv_dumper_1270);
    fifo_csv_dumper_1271 = new("./depth1271.csv");
    cstatus_csv_dumper_1271 = new("./chan_status1271.csv");
    fifo_monitor_1271 = new(fifo_csv_dumper_1271,fifo_intf_1271,cstatus_csv_dumper_1271);
    fifo_csv_dumper_1272 = new("./depth1272.csv");
    cstatus_csv_dumper_1272 = new("./chan_status1272.csv");
    fifo_monitor_1272 = new(fifo_csv_dumper_1272,fifo_intf_1272,cstatus_csv_dumper_1272);
    fifo_csv_dumper_1273 = new("./depth1273.csv");
    cstatus_csv_dumper_1273 = new("./chan_status1273.csv");
    fifo_monitor_1273 = new(fifo_csv_dumper_1273,fifo_intf_1273,cstatus_csv_dumper_1273);
    fifo_csv_dumper_1274 = new("./depth1274.csv");
    cstatus_csv_dumper_1274 = new("./chan_status1274.csv");
    fifo_monitor_1274 = new(fifo_csv_dumper_1274,fifo_intf_1274,cstatus_csv_dumper_1274);
    fifo_csv_dumper_1275 = new("./depth1275.csv");
    cstatus_csv_dumper_1275 = new("./chan_status1275.csv");
    fifo_monitor_1275 = new(fifo_csv_dumper_1275,fifo_intf_1275,cstatus_csv_dumper_1275);
    fifo_csv_dumper_1276 = new("./depth1276.csv");
    cstatus_csv_dumper_1276 = new("./chan_status1276.csv");
    fifo_monitor_1276 = new(fifo_csv_dumper_1276,fifo_intf_1276,cstatus_csv_dumper_1276);
    fifo_csv_dumper_1277 = new("./depth1277.csv");
    cstatus_csv_dumper_1277 = new("./chan_status1277.csv");
    fifo_monitor_1277 = new(fifo_csv_dumper_1277,fifo_intf_1277,cstatus_csv_dumper_1277);
    fifo_csv_dumper_1278 = new("./depth1278.csv");
    cstatus_csv_dumper_1278 = new("./chan_status1278.csv");
    fifo_monitor_1278 = new(fifo_csv_dumper_1278,fifo_intf_1278,cstatus_csv_dumper_1278);
    fifo_csv_dumper_1279 = new("./depth1279.csv");
    cstatus_csv_dumper_1279 = new("./chan_status1279.csv");
    fifo_monitor_1279 = new(fifo_csv_dumper_1279,fifo_intf_1279,cstatus_csv_dumper_1279);
    fifo_csv_dumper_1280 = new("./depth1280.csv");
    cstatus_csv_dumper_1280 = new("./chan_status1280.csv");
    fifo_monitor_1280 = new(fifo_csv_dumper_1280,fifo_intf_1280,cstatus_csv_dumper_1280);
    fifo_csv_dumper_1281 = new("./depth1281.csv");
    cstatus_csv_dumper_1281 = new("./chan_status1281.csv");
    fifo_monitor_1281 = new(fifo_csv_dumper_1281,fifo_intf_1281,cstatus_csv_dumper_1281);
    fifo_csv_dumper_1282 = new("./depth1282.csv");
    cstatus_csv_dumper_1282 = new("./chan_status1282.csv");
    fifo_monitor_1282 = new(fifo_csv_dumper_1282,fifo_intf_1282,cstatus_csv_dumper_1282);
    fifo_csv_dumper_1283 = new("./depth1283.csv");
    cstatus_csv_dumper_1283 = new("./chan_status1283.csv");
    fifo_monitor_1283 = new(fifo_csv_dumper_1283,fifo_intf_1283,cstatus_csv_dumper_1283);
    fifo_csv_dumper_1284 = new("./depth1284.csv");
    cstatus_csv_dumper_1284 = new("./chan_status1284.csv");
    fifo_monitor_1284 = new(fifo_csv_dumper_1284,fifo_intf_1284,cstatus_csv_dumper_1284);
    fifo_csv_dumper_1285 = new("./depth1285.csv");
    cstatus_csv_dumper_1285 = new("./chan_status1285.csv");
    fifo_monitor_1285 = new(fifo_csv_dumper_1285,fifo_intf_1285,cstatus_csv_dumper_1285);
    fifo_csv_dumper_1286 = new("./depth1286.csv");
    cstatus_csv_dumper_1286 = new("./chan_status1286.csv");
    fifo_monitor_1286 = new(fifo_csv_dumper_1286,fifo_intf_1286,cstatus_csv_dumper_1286);
    fifo_csv_dumper_1287 = new("./depth1287.csv");
    cstatus_csv_dumper_1287 = new("./chan_status1287.csv");
    fifo_monitor_1287 = new(fifo_csv_dumper_1287,fifo_intf_1287,cstatus_csv_dumper_1287);
    fifo_csv_dumper_1288 = new("./depth1288.csv");
    cstatus_csv_dumper_1288 = new("./chan_status1288.csv");
    fifo_monitor_1288 = new(fifo_csv_dumper_1288,fifo_intf_1288,cstatus_csv_dumper_1288);
    fifo_csv_dumper_1289 = new("./depth1289.csv");
    cstatus_csv_dumper_1289 = new("./chan_status1289.csv");
    fifo_monitor_1289 = new(fifo_csv_dumper_1289,fifo_intf_1289,cstatus_csv_dumper_1289);
    fifo_csv_dumper_1290 = new("./depth1290.csv");
    cstatus_csv_dumper_1290 = new("./chan_status1290.csv");
    fifo_monitor_1290 = new(fifo_csv_dumper_1290,fifo_intf_1290,cstatus_csv_dumper_1290);
    fifo_csv_dumper_1291 = new("./depth1291.csv");
    cstatus_csv_dumper_1291 = new("./chan_status1291.csv");
    fifo_monitor_1291 = new(fifo_csv_dumper_1291,fifo_intf_1291,cstatus_csv_dumper_1291);
    fifo_csv_dumper_1292 = new("./depth1292.csv");
    cstatus_csv_dumper_1292 = new("./chan_status1292.csv");
    fifo_monitor_1292 = new(fifo_csv_dumper_1292,fifo_intf_1292,cstatus_csv_dumper_1292);
    fifo_csv_dumper_1293 = new("./depth1293.csv");
    cstatus_csv_dumper_1293 = new("./chan_status1293.csv");
    fifo_monitor_1293 = new(fifo_csv_dumper_1293,fifo_intf_1293,cstatus_csv_dumper_1293);
    fifo_csv_dumper_1294 = new("./depth1294.csv");
    cstatus_csv_dumper_1294 = new("./chan_status1294.csv");
    fifo_monitor_1294 = new(fifo_csv_dumper_1294,fifo_intf_1294,cstatus_csv_dumper_1294);
    fifo_csv_dumper_1295 = new("./depth1295.csv");
    cstatus_csv_dumper_1295 = new("./chan_status1295.csv");
    fifo_monitor_1295 = new(fifo_csv_dumper_1295,fifo_intf_1295,cstatus_csv_dumper_1295);
    fifo_csv_dumper_1296 = new("./depth1296.csv");
    cstatus_csv_dumper_1296 = new("./chan_status1296.csv");
    fifo_monitor_1296 = new(fifo_csv_dumper_1296,fifo_intf_1296,cstatus_csv_dumper_1296);
    fifo_csv_dumper_1297 = new("./depth1297.csv");
    cstatus_csv_dumper_1297 = new("./chan_status1297.csv");
    fifo_monitor_1297 = new(fifo_csv_dumper_1297,fifo_intf_1297,cstatus_csv_dumper_1297);
    fifo_csv_dumper_1298 = new("./depth1298.csv");
    cstatus_csv_dumper_1298 = new("./chan_status1298.csv");
    fifo_monitor_1298 = new(fifo_csv_dumper_1298,fifo_intf_1298,cstatus_csv_dumper_1298);
    fifo_csv_dumper_1299 = new("./depth1299.csv");
    cstatus_csv_dumper_1299 = new("./chan_status1299.csv");
    fifo_monitor_1299 = new(fifo_csv_dumper_1299,fifo_intf_1299,cstatus_csv_dumper_1299);
    fifo_csv_dumper_1300 = new("./depth1300.csv");
    cstatus_csv_dumper_1300 = new("./chan_status1300.csv");
    fifo_monitor_1300 = new(fifo_csv_dumper_1300,fifo_intf_1300,cstatus_csv_dumper_1300);
    fifo_csv_dumper_1301 = new("./depth1301.csv");
    cstatus_csv_dumper_1301 = new("./chan_status1301.csv");
    fifo_monitor_1301 = new(fifo_csv_dumper_1301,fifo_intf_1301,cstatus_csv_dumper_1301);
    fifo_csv_dumper_1302 = new("./depth1302.csv");
    cstatus_csv_dumper_1302 = new("./chan_status1302.csv");
    fifo_monitor_1302 = new(fifo_csv_dumper_1302,fifo_intf_1302,cstatus_csv_dumper_1302);
    fifo_csv_dumper_1303 = new("./depth1303.csv");
    cstatus_csv_dumper_1303 = new("./chan_status1303.csv");
    fifo_monitor_1303 = new(fifo_csv_dumper_1303,fifo_intf_1303,cstatus_csv_dumper_1303);
    fifo_csv_dumper_1304 = new("./depth1304.csv");
    cstatus_csv_dumper_1304 = new("./chan_status1304.csv");
    fifo_monitor_1304 = new(fifo_csv_dumper_1304,fifo_intf_1304,cstatus_csv_dumper_1304);
    fifo_csv_dumper_1305 = new("./depth1305.csv");
    cstatus_csv_dumper_1305 = new("./chan_status1305.csv");
    fifo_monitor_1305 = new(fifo_csv_dumper_1305,fifo_intf_1305,cstatus_csv_dumper_1305);
    fifo_csv_dumper_1306 = new("./depth1306.csv");
    cstatus_csv_dumper_1306 = new("./chan_status1306.csv");
    fifo_monitor_1306 = new(fifo_csv_dumper_1306,fifo_intf_1306,cstatus_csv_dumper_1306);
    fifo_csv_dumper_1307 = new("./depth1307.csv");
    cstatus_csv_dumper_1307 = new("./chan_status1307.csv");
    fifo_monitor_1307 = new(fifo_csv_dumper_1307,fifo_intf_1307,cstatus_csv_dumper_1307);
    fifo_csv_dumper_1308 = new("./depth1308.csv");
    cstatus_csv_dumper_1308 = new("./chan_status1308.csv");
    fifo_monitor_1308 = new(fifo_csv_dumper_1308,fifo_intf_1308,cstatus_csv_dumper_1308);
    fifo_csv_dumper_1309 = new("./depth1309.csv");
    cstatus_csv_dumper_1309 = new("./chan_status1309.csv");
    fifo_monitor_1309 = new(fifo_csv_dumper_1309,fifo_intf_1309,cstatus_csv_dumper_1309);
    fifo_csv_dumper_1310 = new("./depth1310.csv");
    cstatus_csv_dumper_1310 = new("./chan_status1310.csv");
    fifo_monitor_1310 = new(fifo_csv_dumper_1310,fifo_intf_1310,cstatus_csv_dumper_1310);
    fifo_csv_dumper_1311 = new("./depth1311.csv");
    cstatus_csv_dumper_1311 = new("./chan_status1311.csv");
    fifo_monitor_1311 = new(fifo_csv_dumper_1311,fifo_intf_1311,cstatus_csv_dumper_1311);
    fifo_csv_dumper_1312 = new("./depth1312.csv");
    cstatus_csv_dumper_1312 = new("./chan_status1312.csv");
    fifo_monitor_1312 = new(fifo_csv_dumper_1312,fifo_intf_1312,cstatus_csv_dumper_1312);
    fifo_csv_dumper_1313 = new("./depth1313.csv");
    cstatus_csv_dumper_1313 = new("./chan_status1313.csv");
    fifo_monitor_1313 = new(fifo_csv_dumper_1313,fifo_intf_1313,cstatus_csv_dumper_1313);
    fifo_csv_dumper_1314 = new("./depth1314.csv");
    cstatus_csv_dumper_1314 = new("./chan_status1314.csv");
    fifo_monitor_1314 = new(fifo_csv_dumper_1314,fifo_intf_1314,cstatus_csv_dumper_1314);
    fifo_csv_dumper_1315 = new("./depth1315.csv");
    cstatus_csv_dumper_1315 = new("./chan_status1315.csv");
    fifo_monitor_1315 = new(fifo_csv_dumper_1315,fifo_intf_1315,cstatus_csv_dumper_1315);
    fifo_csv_dumper_1316 = new("./depth1316.csv");
    cstatus_csv_dumper_1316 = new("./chan_status1316.csv");
    fifo_monitor_1316 = new(fifo_csv_dumper_1316,fifo_intf_1316,cstatus_csv_dumper_1316);
    fifo_csv_dumper_1317 = new("./depth1317.csv");
    cstatus_csv_dumper_1317 = new("./chan_status1317.csv");
    fifo_monitor_1317 = new(fifo_csv_dumper_1317,fifo_intf_1317,cstatus_csv_dumper_1317);
    fifo_csv_dumper_1318 = new("./depth1318.csv");
    cstatus_csv_dumper_1318 = new("./chan_status1318.csv");
    fifo_monitor_1318 = new(fifo_csv_dumper_1318,fifo_intf_1318,cstatus_csv_dumper_1318);
    fifo_csv_dumper_1319 = new("./depth1319.csv");
    cstatus_csv_dumper_1319 = new("./chan_status1319.csv");
    fifo_monitor_1319 = new(fifo_csv_dumper_1319,fifo_intf_1319,cstatus_csv_dumper_1319);
    fifo_csv_dumper_1320 = new("./depth1320.csv");
    cstatus_csv_dumper_1320 = new("./chan_status1320.csv");
    fifo_monitor_1320 = new(fifo_csv_dumper_1320,fifo_intf_1320,cstatus_csv_dumper_1320);
    fifo_csv_dumper_1321 = new("./depth1321.csv");
    cstatus_csv_dumper_1321 = new("./chan_status1321.csv");
    fifo_monitor_1321 = new(fifo_csv_dumper_1321,fifo_intf_1321,cstatus_csv_dumper_1321);
    fifo_csv_dumper_1322 = new("./depth1322.csv");
    cstatus_csv_dumper_1322 = new("./chan_status1322.csv");
    fifo_monitor_1322 = new(fifo_csv_dumper_1322,fifo_intf_1322,cstatus_csv_dumper_1322);
    fifo_csv_dumper_1323 = new("./depth1323.csv");
    cstatus_csv_dumper_1323 = new("./chan_status1323.csv");
    fifo_monitor_1323 = new(fifo_csv_dumper_1323,fifo_intf_1323,cstatus_csv_dumper_1323);
    fifo_csv_dumper_1324 = new("./depth1324.csv");
    cstatus_csv_dumper_1324 = new("./chan_status1324.csv");
    fifo_monitor_1324 = new(fifo_csv_dumper_1324,fifo_intf_1324,cstatus_csv_dumper_1324);
    fifo_csv_dumper_1325 = new("./depth1325.csv");
    cstatus_csv_dumper_1325 = new("./chan_status1325.csv");
    fifo_monitor_1325 = new(fifo_csv_dumper_1325,fifo_intf_1325,cstatus_csv_dumper_1325);
    fifo_csv_dumper_1326 = new("./depth1326.csv");
    cstatus_csv_dumper_1326 = new("./chan_status1326.csv");
    fifo_monitor_1326 = new(fifo_csv_dumper_1326,fifo_intf_1326,cstatus_csv_dumper_1326);
    fifo_csv_dumper_1327 = new("./depth1327.csv");
    cstatus_csv_dumper_1327 = new("./chan_status1327.csv");
    fifo_monitor_1327 = new(fifo_csv_dumper_1327,fifo_intf_1327,cstatus_csv_dumper_1327);
    fifo_csv_dumper_1328 = new("./depth1328.csv");
    cstatus_csv_dumper_1328 = new("./chan_status1328.csv");
    fifo_monitor_1328 = new(fifo_csv_dumper_1328,fifo_intf_1328,cstatus_csv_dumper_1328);
    fifo_csv_dumper_1329 = new("./depth1329.csv");
    cstatus_csv_dumper_1329 = new("./chan_status1329.csv");
    fifo_monitor_1329 = new(fifo_csv_dumper_1329,fifo_intf_1329,cstatus_csv_dumper_1329);
    fifo_csv_dumper_1330 = new("./depth1330.csv");
    cstatus_csv_dumper_1330 = new("./chan_status1330.csv");
    fifo_monitor_1330 = new(fifo_csv_dumper_1330,fifo_intf_1330,cstatus_csv_dumper_1330);
    fifo_csv_dumper_1331 = new("./depth1331.csv");
    cstatus_csv_dumper_1331 = new("./chan_status1331.csv");
    fifo_monitor_1331 = new(fifo_csv_dumper_1331,fifo_intf_1331,cstatus_csv_dumper_1331);
    fifo_csv_dumper_1332 = new("./depth1332.csv");
    cstatus_csv_dumper_1332 = new("./chan_status1332.csv");
    fifo_monitor_1332 = new(fifo_csv_dumper_1332,fifo_intf_1332,cstatus_csv_dumper_1332);
    fifo_csv_dumper_1333 = new("./depth1333.csv");
    cstatus_csv_dumper_1333 = new("./chan_status1333.csv");
    fifo_monitor_1333 = new(fifo_csv_dumper_1333,fifo_intf_1333,cstatus_csv_dumper_1333);
    fifo_csv_dumper_1334 = new("./depth1334.csv");
    cstatus_csv_dumper_1334 = new("./chan_status1334.csv");
    fifo_monitor_1334 = new(fifo_csv_dumper_1334,fifo_intf_1334,cstatus_csv_dumper_1334);
    fifo_csv_dumper_1335 = new("./depth1335.csv");
    cstatus_csv_dumper_1335 = new("./chan_status1335.csv");
    fifo_monitor_1335 = new(fifo_csv_dumper_1335,fifo_intf_1335,cstatus_csv_dumper_1335);
    fifo_csv_dumper_1336 = new("./depth1336.csv");
    cstatus_csv_dumper_1336 = new("./chan_status1336.csv");
    fifo_monitor_1336 = new(fifo_csv_dumper_1336,fifo_intf_1336,cstatus_csv_dumper_1336);
    fifo_csv_dumper_1337 = new("./depth1337.csv");
    cstatus_csv_dumper_1337 = new("./chan_status1337.csv");
    fifo_monitor_1337 = new(fifo_csv_dumper_1337,fifo_intf_1337,cstatus_csv_dumper_1337);
    fifo_csv_dumper_1338 = new("./depth1338.csv");
    cstatus_csv_dumper_1338 = new("./chan_status1338.csv");
    fifo_monitor_1338 = new(fifo_csv_dumper_1338,fifo_intf_1338,cstatus_csv_dumper_1338);
    fifo_csv_dumper_1339 = new("./depth1339.csv");
    cstatus_csv_dumper_1339 = new("./chan_status1339.csv");
    fifo_monitor_1339 = new(fifo_csv_dumper_1339,fifo_intf_1339,cstatus_csv_dumper_1339);
    fifo_csv_dumper_1340 = new("./depth1340.csv");
    cstatus_csv_dumper_1340 = new("./chan_status1340.csv");
    fifo_monitor_1340 = new(fifo_csv_dumper_1340,fifo_intf_1340,cstatus_csv_dumper_1340);
    fifo_csv_dumper_1341 = new("./depth1341.csv");
    cstatus_csv_dumper_1341 = new("./chan_status1341.csv");
    fifo_monitor_1341 = new(fifo_csv_dumper_1341,fifo_intf_1341,cstatus_csv_dumper_1341);
    fifo_csv_dumper_1342 = new("./depth1342.csv");
    cstatus_csv_dumper_1342 = new("./chan_status1342.csv");
    fifo_monitor_1342 = new(fifo_csv_dumper_1342,fifo_intf_1342,cstatus_csv_dumper_1342);
    fifo_csv_dumper_1343 = new("./depth1343.csv");
    cstatus_csv_dumper_1343 = new("./chan_status1343.csv");
    fifo_monitor_1343 = new(fifo_csv_dumper_1343,fifo_intf_1343,cstatus_csv_dumper_1343);
    fifo_csv_dumper_1344 = new("./depth1344.csv");
    cstatus_csv_dumper_1344 = new("./chan_status1344.csv");
    fifo_monitor_1344 = new(fifo_csv_dumper_1344,fifo_intf_1344,cstatus_csv_dumper_1344);
    fifo_csv_dumper_1345 = new("./depth1345.csv");
    cstatus_csv_dumper_1345 = new("./chan_status1345.csv");
    fifo_monitor_1345 = new(fifo_csv_dumper_1345,fifo_intf_1345,cstatus_csv_dumper_1345);
    fifo_csv_dumper_1346 = new("./depth1346.csv");
    cstatus_csv_dumper_1346 = new("./chan_status1346.csv");
    fifo_monitor_1346 = new(fifo_csv_dumper_1346,fifo_intf_1346,cstatus_csv_dumper_1346);
    fifo_csv_dumper_1347 = new("./depth1347.csv");
    cstatus_csv_dumper_1347 = new("./chan_status1347.csv");
    fifo_monitor_1347 = new(fifo_csv_dumper_1347,fifo_intf_1347,cstatus_csv_dumper_1347);
    fifo_csv_dumper_1348 = new("./depth1348.csv");
    cstatus_csv_dumper_1348 = new("./chan_status1348.csv");
    fifo_monitor_1348 = new(fifo_csv_dumper_1348,fifo_intf_1348,cstatus_csv_dumper_1348);
    fifo_csv_dumper_1349 = new("./depth1349.csv");
    cstatus_csv_dumper_1349 = new("./chan_status1349.csv");
    fifo_monitor_1349 = new(fifo_csv_dumper_1349,fifo_intf_1349,cstatus_csv_dumper_1349);
    fifo_csv_dumper_1350 = new("./depth1350.csv");
    cstatus_csv_dumper_1350 = new("./chan_status1350.csv");
    fifo_monitor_1350 = new(fifo_csv_dumper_1350,fifo_intf_1350,cstatus_csv_dumper_1350);
    fifo_csv_dumper_1351 = new("./depth1351.csv");
    cstatus_csv_dumper_1351 = new("./chan_status1351.csv");
    fifo_monitor_1351 = new(fifo_csv_dumper_1351,fifo_intf_1351,cstatus_csv_dumper_1351);
    fifo_csv_dumper_1352 = new("./depth1352.csv");
    cstatus_csv_dumper_1352 = new("./chan_status1352.csv");
    fifo_monitor_1352 = new(fifo_csv_dumper_1352,fifo_intf_1352,cstatus_csv_dumper_1352);
    fifo_csv_dumper_1353 = new("./depth1353.csv");
    cstatus_csv_dumper_1353 = new("./chan_status1353.csv");
    fifo_monitor_1353 = new(fifo_csv_dumper_1353,fifo_intf_1353,cstatus_csv_dumper_1353);
    fifo_csv_dumper_1354 = new("./depth1354.csv");
    cstatus_csv_dumper_1354 = new("./chan_status1354.csv");
    fifo_monitor_1354 = new(fifo_csv_dumper_1354,fifo_intf_1354,cstatus_csv_dumper_1354);
    fifo_csv_dumper_1355 = new("./depth1355.csv");
    cstatus_csv_dumper_1355 = new("./chan_status1355.csv");
    fifo_monitor_1355 = new(fifo_csv_dumper_1355,fifo_intf_1355,cstatus_csv_dumper_1355);
    fifo_csv_dumper_1356 = new("./depth1356.csv");
    cstatus_csv_dumper_1356 = new("./chan_status1356.csv");
    fifo_monitor_1356 = new(fifo_csv_dumper_1356,fifo_intf_1356,cstatus_csv_dumper_1356);
    fifo_csv_dumper_1357 = new("./depth1357.csv");
    cstatus_csv_dumper_1357 = new("./chan_status1357.csv");
    fifo_monitor_1357 = new(fifo_csv_dumper_1357,fifo_intf_1357,cstatus_csv_dumper_1357);
    fifo_csv_dumper_1358 = new("./depth1358.csv");
    cstatus_csv_dumper_1358 = new("./chan_status1358.csv");
    fifo_monitor_1358 = new(fifo_csv_dumper_1358,fifo_intf_1358,cstatus_csv_dumper_1358);
    fifo_csv_dumper_1359 = new("./depth1359.csv");
    cstatus_csv_dumper_1359 = new("./chan_status1359.csv");
    fifo_monitor_1359 = new(fifo_csv_dumper_1359,fifo_intf_1359,cstatus_csv_dumper_1359);
    fifo_csv_dumper_1360 = new("./depth1360.csv");
    cstatus_csv_dumper_1360 = new("./chan_status1360.csv");
    fifo_monitor_1360 = new(fifo_csv_dumper_1360,fifo_intf_1360,cstatus_csv_dumper_1360);
    fifo_csv_dumper_1361 = new("./depth1361.csv");
    cstatus_csv_dumper_1361 = new("./chan_status1361.csv");
    fifo_monitor_1361 = new(fifo_csv_dumper_1361,fifo_intf_1361,cstatus_csv_dumper_1361);
    fifo_csv_dumper_1362 = new("./depth1362.csv");
    cstatus_csv_dumper_1362 = new("./chan_status1362.csv");
    fifo_monitor_1362 = new(fifo_csv_dumper_1362,fifo_intf_1362,cstatus_csv_dumper_1362);
    fifo_csv_dumper_1363 = new("./depth1363.csv");
    cstatus_csv_dumper_1363 = new("./chan_status1363.csv");
    fifo_monitor_1363 = new(fifo_csv_dumper_1363,fifo_intf_1363,cstatus_csv_dumper_1363);
    fifo_csv_dumper_1364 = new("./depth1364.csv");
    cstatus_csv_dumper_1364 = new("./chan_status1364.csv");
    fifo_monitor_1364 = new(fifo_csv_dumper_1364,fifo_intf_1364,cstatus_csv_dumper_1364);
    fifo_csv_dumper_1365 = new("./depth1365.csv");
    cstatus_csv_dumper_1365 = new("./chan_status1365.csv");
    fifo_monitor_1365 = new(fifo_csv_dumper_1365,fifo_intf_1365,cstatus_csv_dumper_1365);
    fifo_csv_dumper_1366 = new("./depth1366.csv");
    cstatus_csv_dumper_1366 = new("./chan_status1366.csv");
    fifo_monitor_1366 = new(fifo_csv_dumper_1366,fifo_intf_1366,cstatus_csv_dumper_1366);
    fifo_csv_dumper_1367 = new("./depth1367.csv");
    cstatus_csv_dumper_1367 = new("./chan_status1367.csv");
    fifo_monitor_1367 = new(fifo_csv_dumper_1367,fifo_intf_1367,cstatus_csv_dumper_1367);
    fifo_csv_dumper_1368 = new("./depth1368.csv");
    cstatus_csv_dumper_1368 = new("./chan_status1368.csv");
    fifo_monitor_1368 = new(fifo_csv_dumper_1368,fifo_intf_1368,cstatus_csv_dumper_1368);
    fifo_csv_dumper_1369 = new("./depth1369.csv");
    cstatus_csv_dumper_1369 = new("./chan_status1369.csv");
    fifo_monitor_1369 = new(fifo_csv_dumper_1369,fifo_intf_1369,cstatus_csv_dumper_1369);
    fifo_csv_dumper_1370 = new("./depth1370.csv");
    cstatus_csv_dumper_1370 = new("./chan_status1370.csv");
    fifo_monitor_1370 = new(fifo_csv_dumper_1370,fifo_intf_1370,cstatus_csv_dumper_1370);
    fifo_csv_dumper_1371 = new("./depth1371.csv");
    cstatus_csv_dumper_1371 = new("./chan_status1371.csv");
    fifo_monitor_1371 = new(fifo_csv_dumper_1371,fifo_intf_1371,cstatus_csv_dumper_1371);
    fifo_csv_dumper_1372 = new("./depth1372.csv");
    cstatus_csv_dumper_1372 = new("./chan_status1372.csv");
    fifo_monitor_1372 = new(fifo_csv_dumper_1372,fifo_intf_1372,cstatus_csv_dumper_1372);
    fifo_csv_dumper_1373 = new("./depth1373.csv");
    cstatus_csv_dumper_1373 = new("./chan_status1373.csv");
    fifo_monitor_1373 = new(fifo_csv_dumper_1373,fifo_intf_1373,cstatus_csv_dumper_1373);
    fifo_csv_dumper_1374 = new("./depth1374.csv");
    cstatus_csv_dumper_1374 = new("./chan_status1374.csv");
    fifo_monitor_1374 = new(fifo_csv_dumper_1374,fifo_intf_1374,cstatus_csv_dumper_1374);
    fifo_csv_dumper_1375 = new("./depth1375.csv");
    cstatus_csv_dumper_1375 = new("./chan_status1375.csv");
    fifo_monitor_1375 = new(fifo_csv_dumper_1375,fifo_intf_1375,cstatus_csv_dumper_1375);
    fifo_csv_dumper_1376 = new("./depth1376.csv");
    cstatus_csv_dumper_1376 = new("./chan_status1376.csv");
    fifo_monitor_1376 = new(fifo_csv_dumper_1376,fifo_intf_1376,cstatus_csv_dumper_1376);
    fifo_csv_dumper_1377 = new("./depth1377.csv");
    cstatus_csv_dumper_1377 = new("./chan_status1377.csv");
    fifo_monitor_1377 = new(fifo_csv_dumper_1377,fifo_intf_1377,cstatus_csv_dumper_1377);
    fifo_csv_dumper_1378 = new("./depth1378.csv");
    cstatus_csv_dumper_1378 = new("./chan_status1378.csv");
    fifo_monitor_1378 = new(fifo_csv_dumper_1378,fifo_intf_1378,cstatus_csv_dumper_1378);
    fifo_csv_dumper_1379 = new("./depth1379.csv");
    cstatus_csv_dumper_1379 = new("./chan_status1379.csv");
    fifo_monitor_1379 = new(fifo_csv_dumper_1379,fifo_intf_1379,cstatus_csv_dumper_1379);
    fifo_csv_dumper_1380 = new("./depth1380.csv");
    cstatus_csv_dumper_1380 = new("./chan_status1380.csv");
    fifo_monitor_1380 = new(fifo_csv_dumper_1380,fifo_intf_1380,cstatus_csv_dumper_1380);
    fifo_csv_dumper_1381 = new("./depth1381.csv");
    cstatus_csv_dumper_1381 = new("./chan_status1381.csv");
    fifo_monitor_1381 = new(fifo_csv_dumper_1381,fifo_intf_1381,cstatus_csv_dumper_1381);
    fifo_csv_dumper_1382 = new("./depth1382.csv");
    cstatus_csv_dumper_1382 = new("./chan_status1382.csv");
    fifo_monitor_1382 = new(fifo_csv_dumper_1382,fifo_intf_1382,cstatus_csv_dumper_1382);
    fifo_csv_dumper_1383 = new("./depth1383.csv");
    cstatus_csv_dumper_1383 = new("./chan_status1383.csv");
    fifo_monitor_1383 = new(fifo_csv_dumper_1383,fifo_intf_1383,cstatus_csv_dumper_1383);
    fifo_csv_dumper_1384 = new("./depth1384.csv");
    cstatus_csv_dumper_1384 = new("./chan_status1384.csv");
    fifo_monitor_1384 = new(fifo_csv_dumper_1384,fifo_intf_1384,cstatus_csv_dumper_1384);
    fifo_csv_dumper_1385 = new("./depth1385.csv");
    cstatus_csv_dumper_1385 = new("./chan_status1385.csv");
    fifo_monitor_1385 = new(fifo_csv_dumper_1385,fifo_intf_1385,cstatus_csv_dumper_1385);
    fifo_csv_dumper_1386 = new("./depth1386.csv");
    cstatus_csv_dumper_1386 = new("./chan_status1386.csv");
    fifo_monitor_1386 = new(fifo_csv_dumper_1386,fifo_intf_1386,cstatus_csv_dumper_1386);
    fifo_csv_dumper_1387 = new("./depth1387.csv");
    cstatus_csv_dumper_1387 = new("./chan_status1387.csv");
    fifo_monitor_1387 = new(fifo_csv_dumper_1387,fifo_intf_1387,cstatus_csv_dumper_1387);
    fifo_csv_dumper_1388 = new("./depth1388.csv");
    cstatus_csv_dumper_1388 = new("./chan_status1388.csv");
    fifo_monitor_1388 = new(fifo_csv_dumper_1388,fifo_intf_1388,cstatus_csv_dumper_1388);
    fifo_csv_dumper_1389 = new("./depth1389.csv");
    cstatus_csv_dumper_1389 = new("./chan_status1389.csv");
    fifo_monitor_1389 = new(fifo_csv_dumper_1389,fifo_intf_1389,cstatus_csv_dumper_1389);
    fifo_csv_dumper_1390 = new("./depth1390.csv");
    cstatus_csv_dumper_1390 = new("./chan_status1390.csv");
    fifo_monitor_1390 = new(fifo_csv_dumper_1390,fifo_intf_1390,cstatus_csv_dumper_1390);
    fifo_csv_dumper_1391 = new("./depth1391.csv");
    cstatus_csv_dumper_1391 = new("./chan_status1391.csv");
    fifo_monitor_1391 = new(fifo_csv_dumper_1391,fifo_intf_1391,cstatus_csv_dumper_1391);
    fifo_csv_dumper_1392 = new("./depth1392.csv");
    cstatus_csv_dumper_1392 = new("./chan_status1392.csv");
    fifo_monitor_1392 = new(fifo_csv_dumper_1392,fifo_intf_1392,cstatus_csv_dumper_1392);
    fifo_csv_dumper_1393 = new("./depth1393.csv");
    cstatus_csv_dumper_1393 = new("./chan_status1393.csv");
    fifo_monitor_1393 = new(fifo_csv_dumper_1393,fifo_intf_1393,cstatus_csv_dumper_1393);
    fifo_csv_dumper_1394 = new("./depth1394.csv");
    cstatus_csv_dumper_1394 = new("./chan_status1394.csv");
    fifo_monitor_1394 = new(fifo_csv_dumper_1394,fifo_intf_1394,cstatus_csv_dumper_1394);
    fifo_csv_dumper_1395 = new("./depth1395.csv");
    cstatus_csv_dumper_1395 = new("./chan_status1395.csv");
    fifo_monitor_1395 = new(fifo_csv_dumper_1395,fifo_intf_1395,cstatus_csv_dumper_1395);
    fifo_csv_dumper_1396 = new("./depth1396.csv");
    cstatus_csv_dumper_1396 = new("./chan_status1396.csv");
    fifo_monitor_1396 = new(fifo_csv_dumper_1396,fifo_intf_1396,cstatus_csv_dumper_1396);
    fifo_csv_dumper_1397 = new("./depth1397.csv");
    cstatus_csv_dumper_1397 = new("./chan_status1397.csv");
    fifo_monitor_1397 = new(fifo_csv_dumper_1397,fifo_intf_1397,cstatus_csv_dumper_1397);
    fifo_csv_dumper_1398 = new("./depth1398.csv");
    cstatus_csv_dumper_1398 = new("./chan_status1398.csv");
    fifo_monitor_1398 = new(fifo_csv_dumper_1398,fifo_intf_1398,cstatus_csv_dumper_1398);
    fifo_csv_dumper_1399 = new("./depth1399.csv");
    cstatus_csv_dumper_1399 = new("./chan_status1399.csv");
    fifo_monitor_1399 = new(fifo_csv_dumper_1399,fifo_intf_1399,cstatus_csv_dumper_1399);
    fifo_csv_dumper_1400 = new("./depth1400.csv");
    cstatus_csv_dumper_1400 = new("./chan_status1400.csv");
    fifo_monitor_1400 = new(fifo_csv_dumper_1400,fifo_intf_1400,cstatus_csv_dumper_1400);
    fifo_csv_dumper_1401 = new("./depth1401.csv");
    cstatus_csv_dumper_1401 = new("./chan_status1401.csv");
    fifo_monitor_1401 = new(fifo_csv_dumper_1401,fifo_intf_1401,cstatus_csv_dumper_1401);
    fifo_csv_dumper_1402 = new("./depth1402.csv");
    cstatus_csv_dumper_1402 = new("./chan_status1402.csv");
    fifo_monitor_1402 = new(fifo_csv_dumper_1402,fifo_intf_1402,cstatus_csv_dumper_1402);
    fifo_csv_dumper_1403 = new("./depth1403.csv");
    cstatus_csv_dumper_1403 = new("./chan_status1403.csv");
    fifo_monitor_1403 = new(fifo_csv_dumper_1403,fifo_intf_1403,cstatus_csv_dumper_1403);
    fifo_csv_dumper_1404 = new("./depth1404.csv");
    cstatus_csv_dumper_1404 = new("./chan_status1404.csv");
    fifo_monitor_1404 = new(fifo_csv_dumper_1404,fifo_intf_1404,cstatus_csv_dumper_1404);
    fifo_csv_dumper_1405 = new("./depth1405.csv");
    cstatus_csv_dumper_1405 = new("./chan_status1405.csv");
    fifo_monitor_1405 = new(fifo_csv_dumper_1405,fifo_intf_1405,cstatus_csv_dumper_1405);
    fifo_csv_dumper_1406 = new("./depth1406.csv");
    cstatus_csv_dumper_1406 = new("./chan_status1406.csv");
    fifo_monitor_1406 = new(fifo_csv_dumper_1406,fifo_intf_1406,cstatus_csv_dumper_1406);
    fifo_csv_dumper_1407 = new("./depth1407.csv");
    cstatus_csv_dumper_1407 = new("./chan_status1407.csv");
    fifo_monitor_1407 = new(fifo_csv_dumper_1407,fifo_intf_1407,cstatus_csv_dumper_1407);
    fifo_csv_dumper_1408 = new("./depth1408.csv");
    cstatus_csv_dumper_1408 = new("./chan_status1408.csv");
    fifo_monitor_1408 = new(fifo_csv_dumper_1408,fifo_intf_1408,cstatus_csv_dumper_1408);
    fifo_csv_dumper_1409 = new("./depth1409.csv");
    cstatus_csv_dumper_1409 = new("./chan_status1409.csv");
    fifo_monitor_1409 = new(fifo_csv_dumper_1409,fifo_intf_1409,cstatus_csv_dumper_1409);
    fifo_csv_dumper_1410 = new("./depth1410.csv");
    cstatus_csv_dumper_1410 = new("./chan_status1410.csv");
    fifo_monitor_1410 = new(fifo_csv_dumper_1410,fifo_intf_1410,cstatus_csv_dumper_1410);
    fifo_csv_dumper_1411 = new("./depth1411.csv");
    cstatus_csv_dumper_1411 = new("./chan_status1411.csv");
    fifo_monitor_1411 = new(fifo_csv_dumper_1411,fifo_intf_1411,cstatus_csv_dumper_1411);
    fifo_csv_dumper_1412 = new("./depth1412.csv");
    cstatus_csv_dumper_1412 = new("./chan_status1412.csv");
    fifo_monitor_1412 = new(fifo_csv_dumper_1412,fifo_intf_1412,cstatus_csv_dumper_1412);
    fifo_csv_dumper_1413 = new("./depth1413.csv");
    cstatus_csv_dumper_1413 = new("./chan_status1413.csv");
    fifo_monitor_1413 = new(fifo_csv_dumper_1413,fifo_intf_1413,cstatus_csv_dumper_1413);
    fifo_csv_dumper_1414 = new("./depth1414.csv");
    cstatus_csv_dumper_1414 = new("./chan_status1414.csv");
    fifo_monitor_1414 = new(fifo_csv_dumper_1414,fifo_intf_1414,cstatus_csv_dumper_1414);
    fifo_csv_dumper_1415 = new("./depth1415.csv");
    cstatus_csv_dumper_1415 = new("./chan_status1415.csv");
    fifo_monitor_1415 = new(fifo_csv_dumper_1415,fifo_intf_1415,cstatus_csv_dumper_1415);
    fifo_csv_dumper_1416 = new("./depth1416.csv");
    cstatus_csv_dumper_1416 = new("./chan_status1416.csv");
    fifo_monitor_1416 = new(fifo_csv_dumper_1416,fifo_intf_1416,cstatus_csv_dumper_1416);
    fifo_csv_dumper_1417 = new("./depth1417.csv");
    cstatus_csv_dumper_1417 = new("./chan_status1417.csv");
    fifo_monitor_1417 = new(fifo_csv_dumper_1417,fifo_intf_1417,cstatus_csv_dumper_1417);
    fifo_csv_dumper_1418 = new("./depth1418.csv");
    cstatus_csv_dumper_1418 = new("./chan_status1418.csv");
    fifo_monitor_1418 = new(fifo_csv_dumper_1418,fifo_intf_1418,cstatus_csv_dumper_1418);
    fifo_csv_dumper_1419 = new("./depth1419.csv");
    cstatus_csv_dumper_1419 = new("./chan_status1419.csv");
    fifo_monitor_1419 = new(fifo_csv_dumper_1419,fifo_intf_1419,cstatus_csv_dumper_1419);
    fifo_csv_dumper_1420 = new("./depth1420.csv");
    cstatus_csv_dumper_1420 = new("./chan_status1420.csv");
    fifo_monitor_1420 = new(fifo_csv_dumper_1420,fifo_intf_1420,cstatus_csv_dumper_1420);
    fifo_csv_dumper_1421 = new("./depth1421.csv");
    cstatus_csv_dumper_1421 = new("./chan_status1421.csv");
    fifo_monitor_1421 = new(fifo_csv_dumper_1421,fifo_intf_1421,cstatus_csv_dumper_1421);
    fifo_csv_dumper_1422 = new("./depth1422.csv");
    cstatus_csv_dumper_1422 = new("./chan_status1422.csv");
    fifo_monitor_1422 = new(fifo_csv_dumper_1422,fifo_intf_1422,cstatus_csv_dumper_1422);
    fifo_csv_dumper_1423 = new("./depth1423.csv");
    cstatus_csv_dumper_1423 = new("./chan_status1423.csv");
    fifo_monitor_1423 = new(fifo_csv_dumper_1423,fifo_intf_1423,cstatus_csv_dumper_1423);
    fifo_csv_dumper_1424 = new("./depth1424.csv");
    cstatus_csv_dumper_1424 = new("./chan_status1424.csv");
    fifo_monitor_1424 = new(fifo_csv_dumper_1424,fifo_intf_1424,cstatus_csv_dumper_1424);
    fifo_csv_dumper_1425 = new("./depth1425.csv");
    cstatus_csv_dumper_1425 = new("./chan_status1425.csv");
    fifo_monitor_1425 = new(fifo_csv_dumper_1425,fifo_intf_1425,cstatus_csv_dumper_1425);
    fifo_csv_dumper_1426 = new("./depth1426.csv");
    cstatus_csv_dumper_1426 = new("./chan_status1426.csv");
    fifo_monitor_1426 = new(fifo_csv_dumper_1426,fifo_intf_1426,cstatus_csv_dumper_1426);
    fifo_csv_dumper_1427 = new("./depth1427.csv");
    cstatus_csv_dumper_1427 = new("./chan_status1427.csv");
    fifo_monitor_1427 = new(fifo_csv_dumper_1427,fifo_intf_1427,cstatus_csv_dumper_1427);
    fifo_csv_dumper_1428 = new("./depth1428.csv");
    cstatus_csv_dumper_1428 = new("./chan_status1428.csv");
    fifo_monitor_1428 = new(fifo_csv_dumper_1428,fifo_intf_1428,cstatus_csv_dumper_1428);
    fifo_csv_dumper_1429 = new("./depth1429.csv");
    cstatus_csv_dumper_1429 = new("./chan_status1429.csv");
    fifo_monitor_1429 = new(fifo_csv_dumper_1429,fifo_intf_1429,cstatus_csv_dumper_1429);
    fifo_csv_dumper_1430 = new("./depth1430.csv");
    cstatus_csv_dumper_1430 = new("./chan_status1430.csv");
    fifo_monitor_1430 = new(fifo_csv_dumper_1430,fifo_intf_1430,cstatus_csv_dumper_1430);
    fifo_csv_dumper_1431 = new("./depth1431.csv");
    cstatus_csv_dumper_1431 = new("./chan_status1431.csv");
    fifo_monitor_1431 = new(fifo_csv_dumper_1431,fifo_intf_1431,cstatus_csv_dumper_1431);
    fifo_csv_dumper_1432 = new("./depth1432.csv");
    cstatus_csv_dumper_1432 = new("./chan_status1432.csv");
    fifo_monitor_1432 = new(fifo_csv_dumper_1432,fifo_intf_1432,cstatus_csv_dumper_1432);
    fifo_csv_dumper_1433 = new("./depth1433.csv");
    cstatus_csv_dumper_1433 = new("./chan_status1433.csv");
    fifo_monitor_1433 = new(fifo_csv_dumper_1433,fifo_intf_1433,cstatus_csv_dumper_1433);
    fifo_csv_dumper_1434 = new("./depth1434.csv");
    cstatus_csv_dumper_1434 = new("./chan_status1434.csv");
    fifo_monitor_1434 = new(fifo_csv_dumper_1434,fifo_intf_1434,cstatus_csv_dumper_1434);
    fifo_csv_dumper_1435 = new("./depth1435.csv");
    cstatus_csv_dumper_1435 = new("./chan_status1435.csv");
    fifo_monitor_1435 = new(fifo_csv_dumper_1435,fifo_intf_1435,cstatus_csv_dumper_1435);
    fifo_csv_dumper_1436 = new("./depth1436.csv");
    cstatus_csv_dumper_1436 = new("./chan_status1436.csv");
    fifo_monitor_1436 = new(fifo_csv_dumper_1436,fifo_intf_1436,cstatus_csv_dumper_1436);
    fifo_csv_dumper_1437 = new("./depth1437.csv");
    cstatus_csv_dumper_1437 = new("./chan_status1437.csv");
    fifo_monitor_1437 = new(fifo_csv_dumper_1437,fifo_intf_1437,cstatus_csv_dumper_1437);
    fifo_csv_dumper_1438 = new("./depth1438.csv");
    cstatus_csv_dumper_1438 = new("./chan_status1438.csv");
    fifo_monitor_1438 = new(fifo_csv_dumper_1438,fifo_intf_1438,cstatus_csv_dumper_1438);
    fifo_csv_dumper_1439 = new("./depth1439.csv");
    cstatus_csv_dumper_1439 = new("./chan_status1439.csv");
    fifo_monitor_1439 = new(fifo_csv_dumper_1439,fifo_intf_1439,cstatus_csv_dumper_1439);
    fifo_csv_dumper_1440 = new("./depth1440.csv");
    cstatus_csv_dumper_1440 = new("./chan_status1440.csv");
    fifo_monitor_1440 = new(fifo_csv_dumper_1440,fifo_intf_1440,cstatus_csv_dumper_1440);
    fifo_csv_dumper_1441 = new("./depth1441.csv");
    cstatus_csv_dumper_1441 = new("./chan_status1441.csv");
    fifo_monitor_1441 = new(fifo_csv_dumper_1441,fifo_intf_1441,cstatus_csv_dumper_1441);
    fifo_csv_dumper_1442 = new("./depth1442.csv");
    cstatus_csv_dumper_1442 = new("./chan_status1442.csv");
    fifo_monitor_1442 = new(fifo_csv_dumper_1442,fifo_intf_1442,cstatus_csv_dumper_1442);
    fifo_csv_dumper_1443 = new("./depth1443.csv");
    cstatus_csv_dumper_1443 = new("./chan_status1443.csv");
    fifo_monitor_1443 = new(fifo_csv_dumper_1443,fifo_intf_1443,cstatus_csv_dumper_1443);
    fifo_csv_dumper_1444 = new("./depth1444.csv");
    cstatus_csv_dumper_1444 = new("./chan_status1444.csv");
    fifo_monitor_1444 = new(fifo_csv_dumper_1444,fifo_intf_1444,cstatus_csv_dumper_1444);
    fifo_csv_dumper_1445 = new("./depth1445.csv");
    cstatus_csv_dumper_1445 = new("./chan_status1445.csv");
    fifo_monitor_1445 = new(fifo_csv_dumper_1445,fifo_intf_1445,cstatus_csv_dumper_1445);
    fifo_csv_dumper_1446 = new("./depth1446.csv");
    cstatus_csv_dumper_1446 = new("./chan_status1446.csv");
    fifo_monitor_1446 = new(fifo_csv_dumper_1446,fifo_intf_1446,cstatus_csv_dumper_1446);
    fifo_csv_dumper_1447 = new("./depth1447.csv");
    cstatus_csv_dumper_1447 = new("./chan_status1447.csv");
    fifo_monitor_1447 = new(fifo_csv_dumper_1447,fifo_intf_1447,cstatus_csv_dumper_1447);
    fifo_csv_dumper_1448 = new("./depth1448.csv");
    cstatus_csv_dumper_1448 = new("./chan_status1448.csv");
    fifo_monitor_1448 = new(fifo_csv_dumper_1448,fifo_intf_1448,cstatus_csv_dumper_1448);
    fifo_csv_dumper_1449 = new("./depth1449.csv");
    cstatus_csv_dumper_1449 = new("./chan_status1449.csv");
    fifo_monitor_1449 = new(fifo_csv_dumper_1449,fifo_intf_1449,cstatus_csv_dumper_1449);
    fifo_csv_dumper_1450 = new("./depth1450.csv");
    cstatus_csv_dumper_1450 = new("./chan_status1450.csv");
    fifo_monitor_1450 = new(fifo_csv_dumper_1450,fifo_intf_1450,cstatus_csv_dumper_1450);
    fifo_csv_dumper_1451 = new("./depth1451.csv");
    cstatus_csv_dumper_1451 = new("./chan_status1451.csv");
    fifo_monitor_1451 = new(fifo_csv_dumper_1451,fifo_intf_1451,cstatus_csv_dumper_1451);
    fifo_csv_dumper_1452 = new("./depth1452.csv");
    cstatus_csv_dumper_1452 = new("./chan_status1452.csv");
    fifo_monitor_1452 = new(fifo_csv_dumper_1452,fifo_intf_1452,cstatus_csv_dumper_1452);
    fifo_csv_dumper_1453 = new("./depth1453.csv");
    cstatus_csv_dumper_1453 = new("./chan_status1453.csv");
    fifo_monitor_1453 = new(fifo_csv_dumper_1453,fifo_intf_1453,cstatus_csv_dumper_1453);
    fifo_csv_dumper_1454 = new("./depth1454.csv");
    cstatus_csv_dumper_1454 = new("./chan_status1454.csv");
    fifo_monitor_1454 = new(fifo_csv_dumper_1454,fifo_intf_1454,cstatus_csv_dumper_1454);
    fifo_csv_dumper_1455 = new("./depth1455.csv");
    cstatus_csv_dumper_1455 = new("./chan_status1455.csv");
    fifo_monitor_1455 = new(fifo_csv_dumper_1455,fifo_intf_1455,cstatus_csv_dumper_1455);
    fifo_csv_dumper_1456 = new("./depth1456.csv");
    cstatus_csv_dumper_1456 = new("./chan_status1456.csv");
    fifo_monitor_1456 = new(fifo_csv_dumper_1456,fifo_intf_1456,cstatus_csv_dumper_1456);
    fifo_csv_dumper_1457 = new("./depth1457.csv");
    cstatus_csv_dumper_1457 = new("./chan_status1457.csv");
    fifo_monitor_1457 = new(fifo_csv_dumper_1457,fifo_intf_1457,cstatus_csv_dumper_1457);
    fifo_csv_dumper_1458 = new("./depth1458.csv");
    cstatus_csv_dumper_1458 = new("./chan_status1458.csv");
    fifo_monitor_1458 = new(fifo_csv_dumper_1458,fifo_intf_1458,cstatus_csv_dumper_1458);
    fifo_csv_dumper_1459 = new("./depth1459.csv");
    cstatus_csv_dumper_1459 = new("./chan_status1459.csv");
    fifo_monitor_1459 = new(fifo_csv_dumper_1459,fifo_intf_1459,cstatus_csv_dumper_1459);
    fifo_csv_dumper_1460 = new("./depth1460.csv");
    cstatus_csv_dumper_1460 = new("./chan_status1460.csv");
    fifo_monitor_1460 = new(fifo_csv_dumper_1460,fifo_intf_1460,cstatus_csv_dumper_1460);
    fifo_csv_dumper_1461 = new("./depth1461.csv");
    cstatus_csv_dumper_1461 = new("./chan_status1461.csv");
    fifo_monitor_1461 = new(fifo_csv_dumper_1461,fifo_intf_1461,cstatus_csv_dumper_1461);
    fifo_csv_dumper_1462 = new("./depth1462.csv");
    cstatus_csv_dumper_1462 = new("./chan_status1462.csv");
    fifo_monitor_1462 = new(fifo_csv_dumper_1462,fifo_intf_1462,cstatus_csv_dumper_1462);
    fifo_csv_dumper_1463 = new("./depth1463.csv");
    cstatus_csv_dumper_1463 = new("./chan_status1463.csv");
    fifo_monitor_1463 = new(fifo_csv_dumper_1463,fifo_intf_1463,cstatus_csv_dumper_1463);
    fifo_csv_dumper_1464 = new("./depth1464.csv");
    cstatus_csv_dumper_1464 = new("./chan_status1464.csv");
    fifo_monitor_1464 = new(fifo_csv_dumper_1464,fifo_intf_1464,cstatus_csv_dumper_1464);
    fifo_csv_dumper_1465 = new("./depth1465.csv");
    cstatus_csv_dumper_1465 = new("./chan_status1465.csv");
    fifo_monitor_1465 = new(fifo_csv_dumper_1465,fifo_intf_1465,cstatus_csv_dumper_1465);
    fifo_csv_dumper_1466 = new("./depth1466.csv");
    cstatus_csv_dumper_1466 = new("./chan_status1466.csv");
    fifo_monitor_1466 = new(fifo_csv_dumper_1466,fifo_intf_1466,cstatus_csv_dumper_1466);
    fifo_csv_dumper_1467 = new("./depth1467.csv");
    cstatus_csv_dumper_1467 = new("./chan_status1467.csv");
    fifo_monitor_1467 = new(fifo_csv_dumper_1467,fifo_intf_1467,cstatus_csv_dumper_1467);
    fifo_csv_dumper_1468 = new("./depth1468.csv");
    cstatus_csv_dumper_1468 = new("./chan_status1468.csv");
    fifo_monitor_1468 = new(fifo_csv_dumper_1468,fifo_intf_1468,cstatus_csv_dumper_1468);
    fifo_csv_dumper_1469 = new("./depth1469.csv");
    cstatus_csv_dumper_1469 = new("./chan_status1469.csv");
    fifo_monitor_1469 = new(fifo_csv_dumper_1469,fifo_intf_1469,cstatus_csv_dumper_1469);
    fifo_csv_dumper_1470 = new("./depth1470.csv");
    cstatus_csv_dumper_1470 = new("./chan_status1470.csv");
    fifo_monitor_1470 = new(fifo_csv_dumper_1470,fifo_intf_1470,cstatus_csv_dumper_1470);
    fifo_csv_dumper_1471 = new("./depth1471.csv");
    cstatus_csv_dumper_1471 = new("./chan_status1471.csv");
    fifo_monitor_1471 = new(fifo_csv_dumper_1471,fifo_intf_1471,cstatus_csv_dumper_1471);
    fifo_csv_dumper_1472 = new("./depth1472.csv");
    cstatus_csv_dumper_1472 = new("./chan_status1472.csv");
    fifo_monitor_1472 = new(fifo_csv_dumper_1472,fifo_intf_1472,cstatus_csv_dumper_1472);
    fifo_csv_dumper_1473 = new("./depth1473.csv");
    cstatus_csv_dumper_1473 = new("./chan_status1473.csv");
    fifo_monitor_1473 = new(fifo_csv_dumper_1473,fifo_intf_1473,cstatus_csv_dumper_1473);
    fifo_csv_dumper_1474 = new("./depth1474.csv");
    cstatus_csv_dumper_1474 = new("./chan_status1474.csv");
    fifo_monitor_1474 = new(fifo_csv_dumper_1474,fifo_intf_1474,cstatus_csv_dumper_1474);
    fifo_csv_dumper_1475 = new("./depth1475.csv");
    cstatus_csv_dumper_1475 = new("./chan_status1475.csv");
    fifo_monitor_1475 = new(fifo_csv_dumper_1475,fifo_intf_1475,cstatus_csv_dumper_1475);
    fifo_csv_dumper_1476 = new("./depth1476.csv");
    cstatus_csv_dumper_1476 = new("./chan_status1476.csv");
    fifo_monitor_1476 = new(fifo_csv_dumper_1476,fifo_intf_1476,cstatus_csv_dumper_1476);
    fifo_csv_dumper_1477 = new("./depth1477.csv");
    cstatus_csv_dumper_1477 = new("./chan_status1477.csv");
    fifo_monitor_1477 = new(fifo_csv_dumper_1477,fifo_intf_1477,cstatus_csv_dumper_1477);
    fifo_csv_dumper_1478 = new("./depth1478.csv");
    cstatus_csv_dumper_1478 = new("./chan_status1478.csv");
    fifo_monitor_1478 = new(fifo_csv_dumper_1478,fifo_intf_1478,cstatus_csv_dumper_1478);
    fifo_csv_dumper_1479 = new("./depth1479.csv");
    cstatus_csv_dumper_1479 = new("./chan_status1479.csv");
    fifo_monitor_1479 = new(fifo_csv_dumper_1479,fifo_intf_1479,cstatus_csv_dumper_1479);
    fifo_csv_dumper_1480 = new("./depth1480.csv");
    cstatus_csv_dumper_1480 = new("./chan_status1480.csv");
    fifo_monitor_1480 = new(fifo_csv_dumper_1480,fifo_intf_1480,cstatus_csv_dumper_1480);
    fifo_csv_dumper_1481 = new("./depth1481.csv");
    cstatus_csv_dumper_1481 = new("./chan_status1481.csv");
    fifo_monitor_1481 = new(fifo_csv_dumper_1481,fifo_intf_1481,cstatus_csv_dumper_1481);
    fifo_csv_dumper_1482 = new("./depth1482.csv");
    cstatus_csv_dumper_1482 = new("./chan_status1482.csv");
    fifo_monitor_1482 = new(fifo_csv_dumper_1482,fifo_intf_1482,cstatus_csv_dumper_1482);
    fifo_csv_dumper_1483 = new("./depth1483.csv");
    cstatus_csv_dumper_1483 = new("./chan_status1483.csv");
    fifo_monitor_1483 = new(fifo_csv_dumper_1483,fifo_intf_1483,cstatus_csv_dumper_1483);
    fifo_csv_dumper_1484 = new("./depth1484.csv");
    cstatus_csv_dumper_1484 = new("./chan_status1484.csv");
    fifo_monitor_1484 = new(fifo_csv_dumper_1484,fifo_intf_1484,cstatus_csv_dumper_1484);
    fifo_csv_dumper_1485 = new("./depth1485.csv");
    cstatus_csv_dumper_1485 = new("./chan_status1485.csv");
    fifo_monitor_1485 = new(fifo_csv_dumper_1485,fifo_intf_1485,cstatus_csv_dumper_1485);
    fifo_csv_dumper_1486 = new("./depth1486.csv");
    cstatus_csv_dumper_1486 = new("./chan_status1486.csv");
    fifo_monitor_1486 = new(fifo_csv_dumper_1486,fifo_intf_1486,cstatus_csv_dumper_1486);
    fifo_csv_dumper_1487 = new("./depth1487.csv");
    cstatus_csv_dumper_1487 = new("./chan_status1487.csv");
    fifo_monitor_1487 = new(fifo_csv_dumper_1487,fifo_intf_1487,cstatus_csv_dumper_1487);
    fifo_csv_dumper_1488 = new("./depth1488.csv");
    cstatus_csv_dumper_1488 = new("./chan_status1488.csv");
    fifo_monitor_1488 = new(fifo_csv_dumper_1488,fifo_intf_1488,cstatus_csv_dumper_1488);
    fifo_csv_dumper_1489 = new("./depth1489.csv");
    cstatus_csv_dumper_1489 = new("./chan_status1489.csv");
    fifo_monitor_1489 = new(fifo_csv_dumper_1489,fifo_intf_1489,cstatus_csv_dumper_1489);
    fifo_csv_dumper_1490 = new("./depth1490.csv");
    cstatus_csv_dumper_1490 = new("./chan_status1490.csv");
    fifo_monitor_1490 = new(fifo_csv_dumper_1490,fifo_intf_1490,cstatus_csv_dumper_1490);
    fifo_csv_dumper_1491 = new("./depth1491.csv");
    cstatus_csv_dumper_1491 = new("./chan_status1491.csv");
    fifo_monitor_1491 = new(fifo_csv_dumper_1491,fifo_intf_1491,cstatus_csv_dumper_1491);
    fifo_csv_dumper_1492 = new("./depth1492.csv");
    cstatus_csv_dumper_1492 = new("./chan_status1492.csv");
    fifo_monitor_1492 = new(fifo_csv_dumper_1492,fifo_intf_1492,cstatus_csv_dumper_1492);
    fifo_csv_dumper_1493 = new("./depth1493.csv");
    cstatus_csv_dumper_1493 = new("./chan_status1493.csv");
    fifo_monitor_1493 = new(fifo_csv_dumper_1493,fifo_intf_1493,cstatus_csv_dumper_1493);
    fifo_csv_dumper_1494 = new("./depth1494.csv");
    cstatus_csv_dumper_1494 = new("./chan_status1494.csv");
    fifo_monitor_1494 = new(fifo_csv_dumper_1494,fifo_intf_1494,cstatus_csv_dumper_1494);
    fifo_csv_dumper_1495 = new("./depth1495.csv");
    cstatus_csv_dumper_1495 = new("./chan_status1495.csv");
    fifo_monitor_1495 = new(fifo_csv_dumper_1495,fifo_intf_1495,cstatus_csv_dumper_1495);
    fifo_csv_dumper_1496 = new("./depth1496.csv");
    cstatus_csv_dumper_1496 = new("./chan_status1496.csv");
    fifo_monitor_1496 = new(fifo_csv_dumper_1496,fifo_intf_1496,cstatus_csv_dumper_1496);
    fifo_csv_dumper_1497 = new("./depth1497.csv");
    cstatus_csv_dumper_1497 = new("./chan_status1497.csv");
    fifo_monitor_1497 = new(fifo_csv_dumper_1497,fifo_intf_1497,cstatus_csv_dumper_1497);
    fifo_csv_dumper_1498 = new("./depth1498.csv");
    cstatus_csv_dumper_1498 = new("./chan_status1498.csv");
    fifo_monitor_1498 = new(fifo_csv_dumper_1498,fifo_intf_1498,cstatus_csv_dumper_1498);
    fifo_csv_dumper_1499 = new("./depth1499.csv");
    cstatus_csv_dumper_1499 = new("./chan_status1499.csv");
    fifo_monitor_1499 = new(fifo_csv_dumper_1499,fifo_intf_1499,cstatus_csv_dumper_1499);
    fifo_csv_dumper_1500 = new("./depth1500.csv");
    cstatus_csv_dumper_1500 = new("./chan_status1500.csv");
    fifo_monitor_1500 = new(fifo_csv_dumper_1500,fifo_intf_1500,cstatus_csv_dumper_1500);
    fifo_csv_dumper_1501 = new("./depth1501.csv");
    cstatus_csv_dumper_1501 = new("./chan_status1501.csv");
    fifo_monitor_1501 = new(fifo_csv_dumper_1501,fifo_intf_1501,cstatus_csv_dumper_1501);
    fifo_csv_dumper_1502 = new("./depth1502.csv");
    cstatus_csv_dumper_1502 = new("./chan_status1502.csv");
    fifo_monitor_1502 = new(fifo_csv_dumper_1502,fifo_intf_1502,cstatus_csv_dumper_1502);
    fifo_csv_dumper_1503 = new("./depth1503.csv");
    cstatus_csv_dumper_1503 = new("./chan_status1503.csv");
    fifo_monitor_1503 = new(fifo_csv_dumper_1503,fifo_intf_1503,cstatus_csv_dumper_1503);
    fifo_csv_dumper_1504 = new("./depth1504.csv");
    cstatus_csv_dumper_1504 = new("./chan_status1504.csv");
    fifo_monitor_1504 = new(fifo_csv_dumper_1504,fifo_intf_1504,cstatus_csv_dumper_1504);
    fifo_csv_dumper_1505 = new("./depth1505.csv");
    cstatus_csv_dumper_1505 = new("./chan_status1505.csv");
    fifo_monitor_1505 = new(fifo_csv_dumper_1505,fifo_intf_1505,cstatus_csv_dumper_1505);
    fifo_csv_dumper_1506 = new("./depth1506.csv");
    cstatus_csv_dumper_1506 = new("./chan_status1506.csv");
    fifo_monitor_1506 = new(fifo_csv_dumper_1506,fifo_intf_1506,cstatus_csv_dumper_1506);
    fifo_csv_dumper_1507 = new("./depth1507.csv");
    cstatus_csv_dumper_1507 = new("./chan_status1507.csv");
    fifo_monitor_1507 = new(fifo_csv_dumper_1507,fifo_intf_1507,cstatus_csv_dumper_1507);
    fifo_csv_dumper_1508 = new("./depth1508.csv");
    cstatus_csv_dumper_1508 = new("./chan_status1508.csv");
    fifo_monitor_1508 = new(fifo_csv_dumper_1508,fifo_intf_1508,cstatus_csv_dumper_1508);
    fifo_csv_dumper_1509 = new("./depth1509.csv");
    cstatus_csv_dumper_1509 = new("./chan_status1509.csv");
    fifo_monitor_1509 = new(fifo_csv_dumper_1509,fifo_intf_1509,cstatus_csv_dumper_1509);
    fifo_csv_dumper_1510 = new("./depth1510.csv");
    cstatus_csv_dumper_1510 = new("./chan_status1510.csv");
    fifo_monitor_1510 = new(fifo_csv_dumper_1510,fifo_intf_1510,cstatus_csv_dumper_1510);
    fifo_csv_dumper_1511 = new("./depth1511.csv");
    cstatus_csv_dumper_1511 = new("./chan_status1511.csv");
    fifo_monitor_1511 = new(fifo_csv_dumper_1511,fifo_intf_1511,cstatus_csv_dumper_1511);
    fifo_csv_dumper_1512 = new("./depth1512.csv");
    cstatus_csv_dumper_1512 = new("./chan_status1512.csv");
    fifo_monitor_1512 = new(fifo_csv_dumper_1512,fifo_intf_1512,cstatus_csv_dumper_1512);
    fifo_csv_dumper_1513 = new("./depth1513.csv");
    cstatus_csv_dumper_1513 = new("./chan_status1513.csv");
    fifo_monitor_1513 = new(fifo_csv_dumper_1513,fifo_intf_1513,cstatus_csv_dumper_1513);
    fifo_csv_dumper_1514 = new("./depth1514.csv");
    cstatus_csv_dumper_1514 = new("./chan_status1514.csv");
    fifo_monitor_1514 = new(fifo_csv_dumper_1514,fifo_intf_1514,cstatus_csv_dumper_1514);
    fifo_csv_dumper_1515 = new("./depth1515.csv");
    cstatus_csv_dumper_1515 = new("./chan_status1515.csv");
    fifo_monitor_1515 = new(fifo_csv_dumper_1515,fifo_intf_1515,cstatus_csv_dumper_1515);
    fifo_csv_dumper_1516 = new("./depth1516.csv");
    cstatus_csv_dumper_1516 = new("./chan_status1516.csv");
    fifo_monitor_1516 = new(fifo_csv_dumper_1516,fifo_intf_1516,cstatus_csv_dumper_1516);
    fifo_csv_dumper_1517 = new("./depth1517.csv");
    cstatus_csv_dumper_1517 = new("./chan_status1517.csv");
    fifo_monitor_1517 = new(fifo_csv_dumper_1517,fifo_intf_1517,cstatus_csv_dumper_1517);
    fifo_csv_dumper_1518 = new("./depth1518.csv");
    cstatus_csv_dumper_1518 = new("./chan_status1518.csv");
    fifo_monitor_1518 = new(fifo_csv_dumper_1518,fifo_intf_1518,cstatus_csv_dumper_1518);
    fifo_csv_dumper_1519 = new("./depth1519.csv");
    cstatus_csv_dumper_1519 = new("./chan_status1519.csv");
    fifo_monitor_1519 = new(fifo_csv_dumper_1519,fifo_intf_1519,cstatus_csv_dumper_1519);
    fifo_csv_dumper_1520 = new("./depth1520.csv");
    cstatus_csv_dumper_1520 = new("./chan_status1520.csv");
    fifo_monitor_1520 = new(fifo_csv_dumper_1520,fifo_intf_1520,cstatus_csv_dumper_1520);
    fifo_csv_dumper_1521 = new("./depth1521.csv");
    cstatus_csv_dumper_1521 = new("./chan_status1521.csv");
    fifo_monitor_1521 = new(fifo_csv_dumper_1521,fifo_intf_1521,cstatus_csv_dumper_1521);
    fifo_csv_dumper_1522 = new("./depth1522.csv");
    cstatus_csv_dumper_1522 = new("./chan_status1522.csv");
    fifo_monitor_1522 = new(fifo_csv_dumper_1522,fifo_intf_1522,cstatus_csv_dumper_1522);
    fifo_csv_dumper_1523 = new("./depth1523.csv");
    cstatus_csv_dumper_1523 = new("./chan_status1523.csv");
    fifo_monitor_1523 = new(fifo_csv_dumper_1523,fifo_intf_1523,cstatus_csv_dumper_1523);
    fifo_csv_dumper_1524 = new("./depth1524.csv");
    cstatus_csv_dumper_1524 = new("./chan_status1524.csv");
    fifo_monitor_1524 = new(fifo_csv_dumper_1524,fifo_intf_1524,cstatus_csv_dumper_1524);
    fifo_csv_dumper_1525 = new("./depth1525.csv");
    cstatus_csv_dumper_1525 = new("./chan_status1525.csv");
    fifo_monitor_1525 = new(fifo_csv_dumper_1525,fifo_intf_1525,cstatus_csv_dumper_1525);
    fifo_csv_dumper_1526 = new("./depth1526.csv");
    cstatus_csv_dumper_1526 = new("./chan_status1526.csv");
    fifo_monitor_1526 = new(fifo_csv_dumper_1526,fifo_intf_1526,cstatus_csv_dumper_1526);
    fifo_csv_dumper_1527 = new("./depth1527.csv");
    cstatus_csv_dumper_1527 = new("./chan_status1527.csv");
    fifo_monitor_1527 = new(fifo_csv_dumper_1527,fifo_intf_1527,cstatus_csv_dumper_1527);
    fifo_csv_dumper_1528 = new("./depth1528.csv");
    cstatus_csv_dumper_1528 = new("./chan_status1528.csv");
    fifo_monitor_1528 = new(fifo_csv_dumper_1528,fifo_intf_1528,cstatus_csv_dumper_1528);
    fifo_csv_dumper_1529 = new("./depth1529.csv");
    cstatus_csv_dumper_1529 = new("./chan_status1529.csv");
    fifo_monitor_1529 = new(fifo_csv_dumper_1529,fifo_intf_1529,cstatus_csv_dumper_1529);
    fifo_csv_dumper_1530 = new("./depth1530.csv");
    cstatus_csv_dumper_1530 = new("./chan_status1530.csv");
    fifo_monitor_1530 = new(fifo_csv_dumper_1530,fifo_intf_1530,cstatus_csv_dumper_1530);
    fifo_csv_dumper_1531 = new("./depth1531.csv");
    cstatus_csv_dumper_1531 = new("./chan_status1531.csv");
    fifo_monitor_1531 = new(fifo_csv_dumper_1531,fifo_intf_1531,cstatus_csv_dumper_1531);
    fifo_csv_dumper_1532 = new("./depth1532.csv");
    cstatus_csv_dumper_1532 = new("./chan_status1532.csv");
    fifo_monitor_1532 = new(fifo_csv_dumper_1532,fifo_intf_1532,cstatus_csv_dumper_1532);
    fifo_csv_dumper_1533 = new("./depth1533.csv");
    cstatus_csv_dumper_1533 = new("./chan_status1533.csv");
    fifo_monitor_1533 = new(fifo_csv_dumper_1533,fifo_intf_1533,cstatus_csv_dumper_1533);
    fifo_csv_dumper_1534 = new("./depth1534.csv");
    cstatus_csv_dumper_1534 = new("./chan_status1534.csv");
    fifo_monitor_1534 = new(fifo_csv_dumper_1534,fifo_intf_1534,cstatus_csv_dumper_1534);
    fifo_csv_dumper_1535 = new("./depth1535.csv");
    cstatus_csv_dumper_1535 = new("./chan_status1535.csv");
    fifo_monitor_1535 = new(fifo_csv_dumper_1535,fifo_intf_1535,cstatus_csv_dumper_1535);
    fifo_csv_dumper_1536 = new("./depth1536.csv");
    cstatus_csv_dumper_1536 = new("./chan_status1536.csv");
    fifo_monitor_1536 = new(fifo_csv_dumper_1536,fifo_intf_1536,cstatus_csv_dumper_1536);
    fifo_csv_dumper_1537 = new("./depth1537.csv");
    cstatus_csv_dumper_1537 = new("./chan_status1537.csv");
    fifo_monitor_1537 = new(fifo_csv_dumper_1537,fifo_intf_1537,cstatus_csv_dumper_1537);
    fifo_csv_dumper_1538 = new("./depth1538.csv");
    cstatus_csv_dumper_1538 = new("./chan_status1538.csv");
    fifo_monitor_1538 = new(fifo_csv_dumper_1538,fifo_intf_1538,cstatus_csv_dumper_1538);
    fifo_csv_dumper_1539 = new("./depth1539.csv");
    cstatus_csv_dumper_1539 = new("./chan_status1539.csv");
    fifo_monitor_1539 = new(fifo_csv_dumper_1539,fifo_intf_1539,cstatus_csv_dumper_1539);
    fifo_csv_dumper_1540 = new("./depth1540.csv");
    cstatus_csv_dumper_1540 = new("./chan_status1540.csv");
    fifo_monitor_1540 = new(fifo_csv_dumper_1540,fifo_intf_1540,cstatus_csv_dumper_1540);
    fifo_csv_dumper_1541 = new("./depth1541.csv");
    cstatus_csv_dumper_1541 = new("./chan_status1541.csv");
    fifo_monitor_1541 = new(fifo_csv_dumper_1541,fifo_intf_1541,cstatus_csv_dumper_1541);
    fifo_csv_dumper_1542 = new("./depth1542.csv");
    cstatus_csv_dumper_1542 = new("./chan_status1542.csv");
    fifo_monitor_1542 = new(fifo_csv_dumper_1542,fifo_intf_1542,cstatus_csv_dumper_1542);
    fifo_csv_dumper_1543 = new("./depth1543.csv");
    cstatus_csv_dumper_1543 = new("./chan_status1543.csv");
    fifo_monitor_1543 = new(fifo_csv_dumper_1543,fifo_intf_1543,cstatus_csv_dumper_1543);
    fifo_csv_dumper_1544 = new("./depth1544.csv");
    cstatus_csv_dumper_1544 = new("./chan_status1544.csv");
    fifo_monitor_1544 = new(fifo_csv_dumper_1544,fifo_intf_1544,cstatus_csv_dumper_1544);
    fifo_csv_dumper_1545 = new("./depth1545.csv");
    cstatus_csv_dumper_1545 = new("./chan_status1545.csv");
    fifo_monitor_1545 = new(fifo_csv_dumper_1545,fifo_intf_1545,cstatus_csv_dumper_1545);
    fifo_csv_dumper_1546 = new("./depth1546.csv");
    cstatus_csv_dumper_1546 = new("./chan_status1546.csv");
    fifo_monitor_1546 = new(fifo_csv_dumper_1546,fifo_intf_1546,cstatus_csv_dumper_1546);
    fifo_csv_dumper_1547 = new("./depth1547.csv");
    cstatus_csv_dumper_1547 = new("./chan_status1547.csv");
    fifo_monitor_1547 = new(fifo_csv_dumper_1547,fifo_intf_1547,cstatus_csv_dumper_1547);
    fifo_csv_dumper_1548 = new("./depth1548.csv");
    cstatus_csv_dumper_1548 = new("./chan_status1548.csv");
    fifo_monitor_1548 = new(fifo_csv_dumper_1548,fifo_intf_1548,cstatus_csv_dumper_1548);
    fifo_csv_dumper_1549 = new("./depth1549.csv");
    cstatus_csv_dumper_1549 = new("./chan_status1549.csv");
    fifo_monitor_1549 = new(fifo_csv_dumper_1549,fifo_intf_1549,cstatus_csv_dumper_1549);
    fifo_csv_dumper_1550 = new("./depth1550.csv");
    cstatus_csv_dumper_1550 = new("./chan_status1550.csv");
    fifo_monitor_1550 = new(fifo_csv_dumper_1550,fifo_intf_1550,cstatus_csv_dumper_1550);
    fifo_csv_dumper_1551 = new("./depth1551.csv");
    cstatus_csv_dumper_1551 = new("./chan_status1551.csv");
    fifo_monitor_1551 = new(fifo_csv_dumper_1551,fifo_intf_1551,cstatus_csv_dumper_1551);
    fifo_csv_dumper_1552 = new("./depth1552.csv");
    cstatus_csv_dumper_1552 = new("./chan_status1552.csv");
    fifo_monitor_1552 = new(fifo_csv_dumper_1552,fifo_intf_1552,cstatus_csv_dumper_1552);
    fifo_csv_dumper_1553 = new("./depth1553.csv");
    cstatus_csv_dumper_1553 = new("./chan_status1553.csv");
    fifo_monitor_1553 = new(fifo_csv_dumper_1553,fifo_intf_1553,cstatus_csv_dumper_1553);
    fifo_csv_dumper_1554 = new("./depth1554.csv");
    cstatus_csv_dumper_1554 = new("./chan_status1554.csv");
    fifo_monitor_1554 = new(fifo_csv_dumper_1554,fifo_intf_1554,cstatus_csv_dumper_1554);
    fifo_csv_dumper_1555 = new("./depth1555.csv");
    cstatus_csv_dumper_1555 = new("./chan_status1555.csv");
    fifo_monitor_1555 = new(fifo_csv_dumper_1555,fifo_intf_1555,cstatus_csv_dumper_1555);
    fifo_csv_dumper_1556 = new("./depth1556.csv");
    cstatus_csv_dumper_1556 = new("./chan_status1556.csv");
    fifo_monitor_1556 = new(fifo_csv_dumper_1556,fifo_intf_1556,cstatus_csv_dumper_1556);
    fifo_csv_dumper_1557 = new("./depth1557.csv");
    cstatus_csv_dumper_1557 = new("./chan_status1557.csv");
    fifo_monitor_1557 = new(fifo_csv_dumper_1557,fifo_intf_1557,cstatus_csv_dumper_1557);
    fifo_csv_dumper_1558 = new("./depth1558.csv");
    cstatus_csv_dumper_1558 = new("./chan_status1558.csv");
    fifo_monitor_1558 = new(fifo_csv_dumper_1558,fifo_intf_1558,cstatus_csv_dumper_1558);
    fifo_csv_dumper_1559 = new("./depth1559.csv");
    cstatus_csv_dumper_1559 = new("./chan_status1559.csv");
    fifo_monitor_1559 = new(fifo_csv_dumper_1559,fifo_intf_1559,cstatus_csv_dumper_1559);
    fifo_csv_dumper_1560 = new("./depth1560.csv");
    cstatus_csv_dumper_1560 = new("./chan_status1560.csv");
    fifo_monitor_1560 = new(fifo_csv_dumper_1560,fifo_intf_1560,cstatus_csv_dumper_1560);
    fifo_csv_dumper_1561 = new("./depth1561.csv");
    cstatus_csv_dumper_1561 = new("./chan_status1561.csv");
    fifo_monitor_1561 = new(fifo_csv_dumper_1561,fifo_intf_1561,cstatus_csv_dumper_1561);
    fifo_csv_dumper_1562 = new("./depth1562.csv");
    cstatus_csv_dumper_1562 = new("./chan_status1562.csv");
    fifo_monitor_1562 = new(fifo_csv_dumper_1562,fifo_intf_1562,cstatus_csv_dumper_1562);
    fifo_csv_dumper_1563 = new("./depth1563.csv");
    cstatus_csv_dumper_1563 = new("./chan_status1563.csv");
    fifo_monitor_1563 = new(fifo_csv_dumper_1563,fifo_intf_1563,cstatus_csv_dumper_1563);
    fifo_csv_dumper_1564 = new("./depth1564.csv");
    cstatus_csv_dumper_1564 = new("./chan_status1564.csv");
    fifo_monitor_1564 = new(fifo_csv_dumper_1564,fifo_intf_1564,cstatus_csv_dumper_1564);
    fifo_csv_dumper_1565 = new("./depth1565.csv");
    cstatus_csv_dumper_1565 = new("./chan_status1565.csv");
    fifo_monitor_1565 = new(fifo_csv_dumper_1565,fifo_intf_1565,cstatus_csv_dumper_1565);
    fifo_csv_dumper_1566 = new("./depth1566.csv");
    cstatus_csv_dumper_1566 = new("./chan_status1566.csv");
    fifo_monitor_1566 = new(fifo_csv_dumper_1566,fifo_intf_1566,cstatus_csv_dumper_1566);
    fifo_csv_dumper_1567 = new("./depth1567.csv");
    cstatus_csv_dumper_1567 = new("./chan_status1567.csv");
    fifo_monitor_1567 = new(fifo_csv_dumper_1567,fifo_intf_1567,cstatus_csv_dumper_1567);
    fifo_csv_dumper_1568 = new("./depth1568.csv");
    cstatus_csv_dumper_1568 = new("./chan_status1568.csv");
    fifo_monitor_1568 = new(fifo_csv_dumper_1568,fifo_intf_1568,cstatus_csv_dumper_1568);
    fifo_csv_dumper_1569 = new("./depth1569.csv");
    cstatus_csv_dumper_1569 = new("./chan_status1569.csv");
    fifo_monitor_1569 = new(fifo_csv_dumper_1569,fifo_intf_1569,cstatus_csv_dumper_1569);
    fifo_csv_dumper_1570 = new("./depth1570.csv");
    cstatus_csv_dumper_1570 = new("./chan_status1570.csv");
    fifo_monitor_1570 = new(fifo_csv_dumper_1570,fifo_intf_1570,cstatus_csv_dumper_1570);
    fifo_csv_dumper_1571 = new("./depth1571.csv");
    cstatus_csv_dumper_1571 = new("./chan_status1571.csv");
    fifo_monitor_1571 = new(fifo_csv_dumper_1571,fifo_intf_1571,cstatus_csv_dumper_1571);
    fifo_csv_dumper_1572 = new("./depth1572.csv");
    cstatus_csv_dumper_1572 = new("./chan_status1572.csv");
    fifo_monitor_1572 = new(fifo_csv_dumper_1572,fifo_intf_1572,cstatus_csv_dumper_1572);
    fifo_csv_dumper_1573 = new("./depth1573.csv");
    cstatus_csv_dumper_1573 = new("./chan_status1573.csv");
    fifo_monitor_1573 = new(fifo_csv_dumper_1573,fifo_intf_1573,cstatus_csv_dumper_1573);
    fifo_csv_dumper_1574 = new("./depth1574.csv");
    cstatus_csv_dumper_1574 = new("./chan_status1574.csv");
    fifo_monitor_1574 = new(fifo_csv_dumper_1574,fifo_intf_1574,cstatus_csv_dumper_1574);
    fifo_csv_dumper_1575 = new("./depth1575.csv");
    cstatus_csv_dumper_1575 = new("./chan_status1575.csv");
    fifo_monitor_1575 = new(fifo_csv_dumper_1575,fifo_intf_1575,cstatus_csv_dumper_1575);
    fifo_csv_dumper_1576 = new("./depth1576.csv");
    cstatus_csv_dumper_1576 = new("./chan_status1576.csv");
    fifo_monitor_1576 = new(fifo_csv_dumper_1576,fifo_intf_1576,cstatus_csv_dumper_1576);
    fifo_csv_dumper_1577 = new("./depth1577.csv");
    cstatus_csv_dumper_1577 = new("./chan_status1577.csv");
    fifo_monitor_1577 = new(fifo_csv_dumper_1577,fifo_intf_1577,cstatus_csv_dumper_1577);
    fifo_csv_dumper_1578 = new("./depth1578.csv");
    cstatus_csv_dumper_1578 = new("./chan_status1578.csv");
    fifo_monitor_1578 = new(fifo_csv_dumper_1578,fifo_intf_1578,cstatus_csv_dumper_1578);
    fifo_csv_dumper_1579 = new("./depth1579.csv");
    cstatus_csv_dumper_1579 = new("./chan_status1579.csv");
    fifo_monitor_1579 = new(fifo_csv_dumper_1579,fifo_intf_1579,cstatus_csv_dumper_1579);
    fifo_csv_dumper_1580 = new("./depth1580.csv");
    cstatus_csv_dumper_1580 = new("./chan_status1580.csv");
    fifo_monitor_1580 = new(fifo_csv_dumper_1580,fifo_intf_1580,cstatus_csv_dumper_1580);
    fifo_csv_dumper_1581 = new("./depth1581.csv");
    cstatus_csv_dumper_1581 = new("./chan_status1581.csv");
    fifo_monitor_1581 = new(fifo_csv_dumper_1581,fifo_intf_1581,cstatus_csv_dumper_1581);
    fifo_csv_dumper_1582 = new("./depth1582.csv");
    cstatus_csv_dumper_1582 = new("./chan_status1582.csv");
    fifo_monitor_1582 = new(fifo_csv_dumper_1582,fifo_intf_1582,cstatus_csv_dumper_1582);
    fifo_csv_dumper_1583 = new("./depth1583.csv");
    cstatus_csv_dumper_1583 = new("./chan_status1583.csv");
    fifo_monitor_1583 = new(fifo_csv_dumper_1583,fifo_intf_1583,cstatus_csv_dumper_1583);
    fifo_csv_dumper_1584 = new("./depth1584.csv");
    cstatus_csv_dumper_1584 = new("./chan_status1584.csv");
    fifo_monitor_1584 = new(fifo_csv_dumper_1584,fifo_intf_1584,cstatus_csv_dumper_1584);
    fifo_csv_dumper_1585 = new("./depth1585.csv");
    cstatus_csv_dumper_1585 = new("./chan_status1585.csv");
    fifo_monitor_1585 = new(fifo_csv_dumper_1585,fifo_intf_1585,cstatus_csv_dumper_1585);
    fifo_csv_dumper_1586 = new("./depth1586.csv");
    cstatus_csv_dumper_1586 = new("./chan_status1586.csv");
    fifo_monitor_1586 = new(fifo_csv_dumper_1586,fifo_intf_1586,cstatus_csv_dumper_1586);
    fifo_csv_dumper_1587 = new("./depth1587.csv");
    cstatus_csv_dumper_1587 = new("./chan_status1587.csv");
    fifo_monitor_1587 = new(fifo_csv_dumper_1587,fifo_intf_1587,cstatus_csv_dumper_1587);
    fifo_csv_dumper_1588 = new("./depth1588.csv");
    cstatus_csv_dumper_1588 = new("./chan_status1588.csv");
    fifo_monitor_1588 = new(fifo_csv_dumper_1588,fifo_intf_1588,cstatus_csv_dumper_1588);
    fifo_csv_dumper_1589 = new("./depth1589.csv");
    cstatus_csv_dumper_1589 = new("./chan_status1589.csv");
    fifo_monitor_1589 = new(fifo_csv_dumper_1589,fifo_intf_1589,cstatus_csv_dumper_1589);
    fifo_csv_dumper_1590 = new("./depth1590.csv");
    cstatus_csv_dumper_1590 = new("./chan_status1590.csv");
    fifo_monitor_1590 = new(fifo_csv_dumper_1590,fifo_intf_1590,cstatus_csv_dumper_1590);
    fifo_csv_dumper_1591 = new("./depth1591.csv");
    cstatus_csv_dumper_1591 = new("./chan_status1591.csv");
    fifo_monitor_1591 = new(fifo_csv_dumper_1591,fifo_intf_1591,cstatus_csv_dumper_1591);
    fifo_csv_dumper_1592 = new("./depth1592.csv");
    cstatus_csv_dumper_1592 = new("./chan_status1592.csv");
    fifo_monitor_1592 = new(fifo_csv_dumper_1592,fifo_intf_1592,cstatus_csv_dumper_1592);
    fifo_csv_dumper_1593 = new("./depth1593.csv");
    cstatus_csv_dumper_1593 = new("./chan_status1593.csv");
    fifo_monitor_1593 = new(fifo_csv_dumper_1593,fifo_intf_1593,cstatus_csv_dumper_1593);
    fifo_csv_dumper_1594 = new("./depth1594.csv");
    cstatus_csv_dumper_1594 = new("./chan_status1594.csv");
    fifo_monitor_1594 = new(fifo_csv_dumper_1594,fifo_intf_1594,cstatus_csv_dumper_1594);
    fifo_csv_dumper_1595 = new("./depth1595.csv");
    cstatus_csv_dumper_1595 = new("./chan_status1595.csv");
    fifo_monitor_1595 = new(fifo_csv_dumper_1595,fifo_intf_1595,cstatus_csv_dumper_1595);
    fifo_csv_dumper_1596 = new("./depth1596.csv");
    cstatus_csv_dumper_1596 = new("./chan_status1596.csv");
    fifo_monitor_1596 = new(fifo_csv_dumper_1596,fifo_intf_1596,cstatus_csv_dumper_1596);
    fifo_csv_dumper_1597 = new("./depth1597.csv");
    cstatus_csv_dumper_1597 = new("./chan_status1597.csv");
    fifo_monitor_1597 = new(fifo_csv_dumper_1597,fifo_intf_1597,cstatus_csv_dumper_1597);
    fifo_csv_dumper_1598 = new("./depth1598.csv");
    cstatus_csv_dumper_1598 = new("./chan_status1598.csv");
    fifo_monitor_1598 = new(fifo_csv_dumper_1598,fifo_intf_1598,cstatus_csv_dumper_1598);
    fifo_csv_dumper_1599 = new("./depth1599.csv");
    cstatus_csv_dumper_1599 = new("./chan_status1599.csv");
    fifo_monitor_1599 = new(fifo_csv_dumper_1599,fifo_intf_1599,cstatus_csv_dumper_1599);
    fifo_csv_dumper_1600 = new("./depth1600.csv");
    cstatus_csv_dumper_1600 = new("./chan_status1600.csv");
    fifo_monitor_1600 = new(fifo_csv_dumper_1600,fifo_intf_1600,cstatus_csv_dumper_1600);
    fifo_csv_dumper_1601 = new("./depth1601.csv");
    cstatus_csv_dumper_1601 = new("./chan_status1601.csv");
    fifo_monitor_1601 = new(fifo_csv_dumper_1601,fifo_intf_1601,cstatus_csv_dumper_1601);
    fifo_csv_dumper_1602 = new("./depth1602.csv");
    cstatus_csv_dumper_1602 = new("./chan_status1602.csv");
    fifo_monitor_1602 = new(fifo_csv_dumper_1602,fifo_intf_1602,cstatus_csv_dumper_1602);
    fifo_csv_dumper_1603 = new("./depth1603.csv");
    cstatus_csv_dumper_1603 = new("./chan_status1603.csv");
    fifo_monitor_1603 = new(fifo_csv_dumper_1603,fifo_intf_1603,cstatus_csv_dumper_1603);
    fifo_csv_dumper_1604 = new("./depth1604.csv");
    cstatus_csv_dumper_1604 = new("./chan_status1604.csv");
    fifo_monitor_1604 = new(fifo_csv_dumper_1604,fifo_intf_1604,cstatus_csv_dumper_1604);
    fifo_csv_dumper_1605 = new("./depth1605.csv");
    cstatus_csv_dumper_1605 = new("./chan_status1605.csv");
    fifo_monitor_1605 = new(fifo_csv_dumper_1605,fifo_intf_1605,cstatus_csv_dumper_1605);
    fifo_csv_dumper_1606 = new("./depth1606.csv");
    cstatus_csv_dumper_1606 = new("./chan_status1606.csv");
    fifo_monitor_1606 = new(fifo_csv_dumper_1606,fifo_intf_1606,cstatus_csv_dumper_1606);
    fifo_csv_dumper_1607 = new("./depth1607.csv");
    cstatus_csv_dumper_1607 = new("./chan_status1607.csv");
    fifo_monitor_1607 = new(fifo_csv_dumper_1607,fifo_intf_1607,cstatus_csv_dumper_1607);
    fifo_csv_dumper_1608 = new("./depth1608.csv");
    cstatus_csv_dumper_1608 = new("./chan_status1608.csv");
    fifo_monitor_1608 = new(fifo_csv_dumper_1608,fifo_intf_1608,cstatus_csv_dumper_1608);
    fifo_csv_dumper_1609 = new("./depth1609.csv");
    cstatus_csv_dumper_1609 = new("./chan_status1609.csv");
    fifo_monitor_1609 = new(fifo_csv_dumper_1609,fifo_intf_1609,cstatus_csv_dumper_1609);
    fifo_csv_dumper_1610 = new("./depth1610.csv");
    cstatus_csv_dumper_1610 = new("./chan_status1610.csv");
    fifo_monitor_1610 = new(fifo_csv_dumper_1610,fifo_intf_1610,cstatus_csv_dumper_1610);
    fifo_csv_dumper_1611 = new("./depth1611.csv");
    cstatus_csv_dumper_1611 = new("./chan_status1611.csv");
    fifo_monitor_1611 = new(fifo_csv_dumper_1611,fifo_intf_1611,cstatus_csv_dumper_1611);
    fifo_csv_dumper_1612 = new("./depth1612.csv");
    cstatus_csv_dumper_1612 = new("./chan_status1612.csv");
    fifo_monitor_1612 = new(fifo_csv_dumper_1612,fifo_intf_1612,cstatus_csv_dumper_1612);
    fifo_csv_dumper_1613 = new("./depth1613.csv");
    cstatus_csv_dumper_1613 = new("./chan_status1613.csv");
    fifo_monitor_1613 = new(fifo_csv_dumper_1613,fifo_intf_1613,cstatus_csv_dumper_1613);
    fifo_csv_dumper_1614 = new("./depth1614.csv");
    cstatus_csv_dumper_1614 = new("./chan_status1614.csv");
    fifo_monitor_1614 = new(fifo_csv_dumper_1614,fifo_intf_1614,cstatus_csv_dumper_1614);
    fifo_csv_dumper_1615 = new("./depth1615.csv");
    cstatus_csv_dumper_1615 = new("./chan_status1615.csv");
    fifo_monitor_1615 = new(fifo_csv_dumper_1615,fifo_intf_1615,cstatus_csv_dumper_1615);
    fifo_csv_dumper_1616 = new("./depth1616.csv");
    cstatus_csv_dumper_1616 = new("./chan_status1616.csv");
    fifo_monitor_1616 = new(fifo_csv_dumper_1616,fifo_intf_1616,cstatus_csv_dumper_1616);
    fifo_csv_dumper_1617 = new("./depth1617.csv");
    cstatus_csv_dumper_1617 = new("./chan_status1617.csv");
    fifo_monitor_1617 = new(fifo_csv_dumper_1617,fifo_intf_1617,cstatus_csv_dumper_1617);
    fifo_csv_dumper_1618 = new("./depth1618.csv");
    cstatus_csv_dumper_1618 = new("./chan_status1618.csv");
    fifo_monitor_1618 = new(fifo_csv_dumper_1618,fifo_intf_1618,cstatus_csv_dumper_1618);
    fifo_csv_dumper_1619 = new("./depth1619.csv");
    cstatus_csv_dumper_1619 = new("./chan_status1619.csv");
    fifo_monitor_1619 = new(fifo_csv_dumper_1619,fifo_intf_1619,cstatus_csv_dumper_1619);
    fifo_csv_dumper_1620 = new("./depth1620.csv");
    cstatus_csv_dumper_1620 = new("./chan_status1620.csv");
    fifo_monitor_1620 = new(fifo_csv_dumper_1620,fifo_intf_1620,cstatus_csv_dumper_1620);
    fifo_csv_dumper_1621 = new("./depth1621.csv");
    cstatus_csv_dumper_1621 = new("./chan_status1621.csv");
    fifo_monitor_1621 = new(fifo_csv_dumper_1621,fifo_intf_1621,cstatus_csv_dumper_1621);
    fifo_csv_dumper_1622 = new("./depth1622.csv");
    cstatus_csv_dumper_1622 = new("./chan_status1622.csv");
    fifo_monitor_1622 = new(fifo_csv_dumper_1622,fifo_intf_1622,cstatus_csv_dumper_1622);
    fifo_csv_dumper_1623 = new("./depth1623.csv");
    cstatus_csv_dumper_1623 = new("./chan_status1623.csv");
    fifo_monitor_1623 = new(fifo_csv_dumper_1623,fifo_intf_1623,cstatus_csv_dumper_1623);
    fifo_csv_dumper_1624 = new("./depth1624.csv");
    cstatus_csv_dumper_1624 = new("./chan_status1624.csv");
    fifo_monitor_1624 = new(fifo_csv_dumper_1624,fifo_intf_1624,cstatus_csv_dumper_1624);
    fifo_csv_dumper_1625 = new("./depth1625.csv");
    cstatus_csv_dumper_1625 = new("./chan_status1625.csv");
    fifo_monitor_1625 = new(fifo_csv_dumper_1625,fifo_intf_1625,cstatus_csv_dumper_1625);
    fifo_csv_dumper_1626 = new("./depth1626.csv");
    cstatus_csv_dumper_1626 = new("./chan_status1626.csv");
    fifo_monitor_1626 = new(fifo_csv_dumper_1626,fifo_intf_1626,cstatus_csv_dumper_1626);
    fifo_csv_dumper_1627 = new("./depth1627.csv");
    cstatus_csv_dumper_1627 = new("./chan_status1627.csv");
    fifo_monitor_1627 = new(fifo_csv_dumper_1627,fifo_intf_1627,cstatus_csv_dumper_1627);
    fifo_csv_dumper_1628 = new("./depth1628.csv");
    cstatus_csv_dumper_1628 = new("./chan_status1628.csv");
    fifo_monitor_1628 = new(fifo_csv_dumper_1628,fifo_intf_1628,cstatus_csv_dumper_1628);
    fifo_csv_dumper_1629 = new("./depth1629.csv");
    cstatus_csv_dumper_1629 = new("./chan_status1629.csv");
    fifo_monitor_1629 = new(fifo_csv_dumper_1629,fifo_intf_1629,cstatus_csv_dumper_1629);
    fifo_csv_dumper_1630 = new("./depth1630.csv");
    cstatus_csv_dumper_1630 = new("./chan_status1630.csv");
    fifo_monitor_1630 = new(fifo_csv_dumper_1630,fifo_intf_1630,cstatus_csv_dumper_1630);
    fifo_csv_dumper_1631 = new("./depth1631.csv");
    cstatus_csv_dumper_1631 = new("./chan_status1631.csv");
    fifo_monitor_1631 = new(fifo_csv_dumper_1631,fifo_intf_1631,cstatus_csv_dumper_1631);
    fifo_csv_dumper_1632 = new("./depth1632.csv");
    cstatus_csv_dumper_1632 = new("./chan_status1632.csv");
    fifo_monitor_1632 = new(fifo_csv_dumper_1632,fifo_intf_1632,cstatus_csv_dumper_1632);
    fifo_csv_dumper_1633 = new("./depth1633.csv");
    cstatus_csv_dumper_1633 = new("./chan_status1633.csv");
    fifo_monitor_1633 = new(fifo_csv_dumper_1633,fifo_intf_1633,cstatus_csv_dumper_1633);
    fifo_csv_dumper_1634 = new("./depth1634.csv");
    cstatus_csv_dumper_1634 = new("./chan_status1634.csv");
    fifo_monitor_1634 = new(fifo_csv_dumper_1634,fifo_intf_1634,cstatus_csv_dumper_1634);
    fifo_csv_dumper_1635 = new("./depth1635.csv");
    cstatus_csv_dumper_1635 = new("./chan_status1635.csv");
    fifo_monitor_1635 = new(fifo_csv_dumper_1635,fifo_intf_1635,cstatus_csv_dumper_1635);
    fifo_csv_dumper_1636 = new("./depth1636.csv");
    cstatus_csv_dumper_1636 = new("./chan_status1636.csv");
    fifo_monitor_1636 = new(fifo_csv_dumper_1636,fifo_intf_1636,cstatus_csv_dumper_1636);
    fifo_csv_dumper_1637 = new("./depth1637.csv");
    cstatus_csv_dumper_1637 = new("./chan_status1637.csv");
    fifo_monitor_1637 = new(fifo_csv_dumper_1637,fifo_intf_1637,cstatus_csv_dumper_1637);
    fifo_csv_dumper_1638 = new("./depth1638.csv");
    cstatus_csv_dumper_1638 = new("./chan_status1638.csv");
    fifo_monitor_1638 = new(fifo_csv_dumper_1638,fifo_intf_1638,cstatus_csv_dumper_1638);
    fifo_csv_dumper_1639 = new("./depth1639.csv");
    cstatus_csv_dumper_1639 = new("./chan_status1639.csv");
    fifo_monitor_1639 = new(fifo_csv_dumper_1639,fifo_intf_1639,cstatus_csv_dumper_1639);
    fifo_csv_dumper_1640 = new("./depth1640.csv");
    cstatus_csv_dumper_1640 = new("./chan_status1640.csv");
    fifo_monitor_1640 = new(fifo_csv_dumper_1640,fifo_intf_1640,cstatus_csv_dumper_1640);
    fifo_csv_dumper_1641 = new("./depth1641.csv");
    cstatus_csv_dumper_1641 = new("./chan_status1641.csv");
    fifo_monitor_1641 = new(fifo_csv_dumper_1641,fifo_intf_1641,cstatus_csv_dumper_1641);
    fifo_csv_dumper_1642 = new("./depth1642.csv");
    cstatus_csv_dumper_1642 = new("./chan_status1642.csv");
    fifo_monitor_1642 = new(fifo_csv_dumper_1642,fifo_intf_1642,cstatus_csv_dumper_1642);
    fifo_csv_dumper_1643 = new("./depth1643.csv");
    cstatus_csv_dumper_1643 = new("./chan_status1643.csv");
    fifo_monitor_1643 = new(fifo_csv_dumper_1643,fifo_intf_1643,cstatus_csv_dumper_1643);
    fifo_csv_dumper_1644 = new("./depth1644.csv");
    cstatus_csv_dumper_1644 = new("./chan_status1644.csv");
    fifo_monitor_1644 = new(fifo_csv_dumper_1644,fifo_intf_1644,cstatus_csv_dumper_1644);
    fifo_csv_dumper_1645 = new("./depth1645.csv");
    cstatus_csv_dumper_1645 = new("./chan_status1645.csv");
    fifo_monitor_1645 = new(fifo_csv_dumper_1645,fifo_intf_1645,cstatus_csv_dumper_1645);
    fifo_csv_dumper_1646 = new("./depth1646.csv");
    cstatus_csv_dumper_1646 = new("./chan_status1646.csv");
    fifo_monitor_1646 = new(fifo_csv_dumper_1646,fifo_intf_1646,cstatus_csv_dumper_1646);
    fifo_csv_dumper_1647 = new("./depth1647.csv");
    cstatus_csv_dumper_1647 = new("./chan_status1647.csv");
    fifo_monitor_1647 = new(fifo_csv_dumper_1647,fifo_intf_1647,cstatus_csv_dumper_1647);
    fifo_csv_dumper_1648 = new("./depth1648.csv");
    cstatus_csv_dumper_1648 = new("./chan_status1648.csv");
    fifo_monitor_1648 = new(fifo_csv_dumper_1648,fifo_intf_1648,cstatus_csv_dumper_1648);
    fifo_csv_dumper_1649 = new("./depth1649.csv");
    cstatus_csv_dumper_1649 = new("./chan_status1649.csv");
    fifo_monitor_1649 = new(fifo_csv_dumper_1649,fifo_intf_1649,cstatus_csv_dumper_1649);
    fifo_csv_dumper_1650 = new("./depth1650.csv");
    cstatus_csv_dumper_1650 = new("./chan_status1650.csv");
    fifo_monitor_1650 = new(fifo_csv_dumper_1650,fifo_intf_1650,cstatus_csv_dumper_1650);
    fifo_csv_dumper_1651 = new("./depth1651.csv");
    cstatus_csv_dumper_1651 = new("./chan_status1651.csv");
    fifo_monitor_1651 = new(fifo_csv_dumper_1651,fifo_intf_1651,cstatus_csv_dumper_1651);
    fifo_csv_dumper_1652 = new("./depth1652.csv");
    cstatus_csv_dumper_1652 = new("./chan_status1652.csv");
    fifo_monitor_1652 = new(fifo_csv_dumper_1652,fifo_intf_1652,cstatus_csv_dumper_1652);
    fifo_csv_dumper_1653 = new("./depth1653.csv");
    cstatus_csv_dumper_1653 = new("./chan_status1653.csv");
    fifo_monitor_1653 = new(fifo_csv_dumper_1653,fifo_intf_1653,cstatus_csv_dumper_1653);
    fifo_csv_dumper_1654 = new("./depth1654.csv");
    cstatus_csv_dumper_1654 = new("./chan_status1654.csv");
    fifo_monitor_1654 = new(fifo_csv_dumper_1654,fifo_intf_1654,cstatus_csv_dumper_1654);
    fifo_csv_dumper_1655 = new("./depth1655.csv");
    cstatus_csv_dumper_1655 = new("./chan_status1655.csv");
    fifo_monitor_1655 = new(fifo_csv_dumper_1655,fifo_intf_1655,cstatus_csv_dumper_1655);
    fifo_csv_dumper_1656 = new("./depth1656.csv");
    cstatus_csv_dumper_1656 = new("./chan_status1656.csv");
    fifo_monitor_1656 = new(fifo_csv_dumper_1656,fifo_intf_1656,cstatus_csv_dumper_1656);
    fifo_csv_dumper_1657 = new("./depth1657.csv");
    cstatus_csv_dumper_1657 = new("./chan_status1657.csv");
    fifo_monitor_1657 = new(fifo_csv_dumper_1657,fifo_intf_1657,cstatus_csv_dumper_1657);
    fifo_csv_dumper_1658 = new("./depth1658.csv");
    cstatus_csv_dumper_1658 = new("./chan_status1658.csv");
    fifo_monitor_1658 = new(fifo_csv_dumper_1658,fifo_intf_1658,cstatus_csv_dumper_1658);
    fifo_csv_dumper_1659 = new("./depth1659.csv");
    cstatus_csv_dumper_1659 = new("./chan_status1659.csv");
    fifo_monitor_1659 = new(fifo_csv_dumper_1659,fifo_intf_1659,cstatus_csv_dumper_1659);
    fifo_csv_dumper_1660 = new("./depth1660.csv");
    cstatus_csv_dumper_1660 = new("./chan_status1660.csv");
    fifo_monitor_1660 = new(fifo_csv_dumper_1660,fifo_intf_1660,cstatus_csv_dumper_1660);
    fifo_csv_dumper_1661 = new("./depth1661.csv");
    cstatus_csv_dumper_1661 = new("./chan_status1661.csv");
    fifo_monitor_1661 = new(fifo_csv_dumper_1661,fifo_intf_1661,cstatus_csv_dumper_1661);
    fifo_csv_dumper_1662 = new("./depth1662.csv");
    cstatus_csv_dumper_1662 = new("./chan_status1662.csv");
    fifo_monitor_1662 = new(fifo_csv_dumper_1662,fifo_intf_1662,cstatus_csv_dumper_1662);
    fifo_csv_dumper_1663 = new("./depth1663.csv");
    cstatus_csv_dumper_1663 = new("./chan_status1663.csv");
    fifo_monitor_1663 = new(fifo_csv_dumper_1663,fifo_intf_1663,cstatus_csv_dumper_1663);
    fifo_csv_dumper_1664 = new("./depth1664.csv");
    cstatus_csv_dumper_1664 = new("./chan_status1664.csv");
    fifo_monitor_1664 = new(fifo_csv_dumper_1664,fifo_intf_1664,cstatus_csv_dumper_1664);
    fifo_csv_dumper_1665 = new("./depth1665.csv");
    cstatus_csv_dumper_1665 = new("./chan_status1665.csv");
    fifo_monitor_1665 = new(fifo_csv_dumper_1665,fifo_intf_1665,cstatus_csv_dumper_1665);
    fifo_csv_dumper_1666 = new("./depth1666.csv");
    cstatus_csv_dumper_1666 = new("./chan_status1666.csv");
    fifo_monitor_1666 = new(fifo_csv_dumper_1666,fifo_intf_1666,cstatus_csv_dumper_1666);
    fifo_csv_dumper_1667 = new("./depth1667.csv");
    cstatus_csv_dumper_1667 = new("./chan_status1667.csv");
    fifo_monitor_1667 = new(fifo_csv_dumper_1667,fifo_intf_1667,cstatus_csv_dumper_1667);
    fifo_csv_dumper_1668 = new("./depth1668.csv");
    cstatus_csv_dumper_1668 = new("./chan_status1668.csv");
    fifo_monitor_1668 = new(fifo_csv_dumper_1668,fifo_intf_1668,cstatus_csv_dumper_1668);
    fifo_csv_dumper_1669 = new("./depth1669.csv");
    cstatus_csv_dumper_1669 = new("./chan_status1669.csv");
    fifo_monitor_1669 = new(fifo_csv_dumper_1669,fifo_intf_1669,cstatus_csv_dumper_1669);
    fifo_csv_dumper_1670 = new("./depth1670.csv");
    cstatus_csv_dumper_1670 = new("./chan_status1670.csv");
    fifo_monitor_1670 = new(fifo_csv_dumper_1670,fifo_intf_1670,cstatus_csv_dumper_1670);
    fifo_csv_dumper_1671 = new("./depth1671.csv");
    cstatus_csv_dumper_1671 = new("./chan_status1671.csv");
    fifo_monitor_1671 = new(fifo_csv_dumper_1671,fifo_intf_1671,cstatus_csv_dumper_1671);
    fifo_csv_dumper_1672 = new("./depth1672.csv");
    cstatus_csv_dumper_1672 = new("./chan_status1672.csv");
    fifo_monitor_1672 = new(fifo_csv_dumper_1672,fifo_intf_1672,cstatus_csv_dumper_1672);
    fifo_csv_dumper_1673 = new("./depth1673.csv");
    cstatus_csv_dumper_1673 = new("./chan_status1673.csv");
    fifo_monitor_1673 = new(fifo_csv_dumper_1673,fifo_intf_1673,cstatus_csv_dumper_1673);
    fifo_csv_dumper_1674 = new("./depth1674.csv");
    cstatus_csv_dumper_1674 = new("./chan_status1674.csv");
    fifo_monitor_1674 = new(fifo_csv_dumper_1674,fifo_intf_1674,cstatus_csv_dumper_1674);
    fifo_csv_dumper_1675 = new("./depth1675.csv");
    cstatus_csv_dumper_1675 = new("./chan_status1675.csv");
    fifo_monitor_1675 = new(fifo_csv_dumper_1675,fifo_intf_1675,cstatus_csv_dumper_1675);
    fifo_csv_dumper_1676 = new("./depth1676.csv");
    cstatus_csv_dumper_1676 = new("./chan_status1676.csv");
    fifo_monitor_1676 = new(fifo_csv_dumper_1676,fifo_intf_1676,cstatus_csv_dumper_1676);
    fifo_csv_dumper_1677 = new("./depth1677.csv");
    cstatus_csv_dumper_1677 = new("./chan_status1677.csv");
    fifo_monitor_1677 = new(fifo_csv_dumper_1677,fifo_intf_1677,cstatus_csv_dumper_1677);
    fifo_csv_dumper_1678 = new("./depth1678.csv");
    cstatus_csv_dumper_1678 = new("./chan_status1678.csv");
    fifo_monitor_1678 = new(fifo_csv_dumper_1678,fifo_intf_1678,cstatus_csv_dumper_1678);
    fifo_csv_dumper_1679 = new("./depth1679.csv");
    cstatus_csv_dumper_1679 = new("./chan_status1679.csv");
    fifo_monitor_1679 = new(fifo_csv_dumper_1679,fifo_intf_1679,cstatus_csv_dumper_1679);
    fifo_csv_dumper_1680 = new("./depth1680.csv");
    cstatus_csv_dumper_1680 = new("./chan_status1680.csv");
    fifo_monitor_1680 = new(fifo_csv_dumper_1680,fifo_intf_1680,cstatus_csv_dumper_1680);
    fifo_csv_dumper_1681 = new("./depth1681.csv");
    cstatus_csv_dumper_1681 = new("./chan_status1681.csv");
    fifo_monitor_1681 = new(fifo_csv_dumper_1681,fifo_intf_1681,cstatus_csv_dumper_1681);
    fifo_csv_dumper_1682 = new("./depth1682.csv");
    cstatus_csv_dumper_1682 = new("./chan_status1682.csv");
    fifo_monitor_1682 = new(fifo_csv_dumper_1682,fifo_intf_1682,cstatus_csv_dumper_1682);
    fifo_csv_dumper_1683 = new("./depth1683.csv");
    cstatus_csv_dumper_1683 = new("./chan_status1683.csv");
    fifo_monitor_1683 = new(fifo_csv_dumper_1683,fifo_intf_1683,cstatus_csv_dumper_1683);
    fifo_csv_dumper_1684 = new("./depth1684.csv");
    cstatus_csv_dumper_1684 = new("./chan_status1684.csv");
    fifo_monitor_1684 = new(fifo_csv_dumper_1684,fifo_intf_1684,cstatus_csv_dumper_1684);
    fifo_csv_dumper_1685 = new("./depth1685.csv");
    cstatus_csv_dumper_1685 = new("./chan_status1685.csv");
    fifo_monitor_1685 = new(fifo_csv_dumper_1685,fifo_intf_1685,cstatus_csv_dumper_1685);
    fifo_csv_dumper_1686 = new("./depth1686.csv");
    cstatus_csv_dumper_1686 = new("./chan_status1686.csv");
    fifo_monitor_1686 = new(fifo_csv_dumper_1686,fifo_intf_1686,cstatus_csv_dumper_1686);
    fifo_csv_dumper_1687 = new("./depth1687.csv");
    cstatus_csv_dumper_1687 = new("./chan_status1687.csv");
    fifo_monitor_1687 = new(fifo_csv_dumper_1687,fifo_intf_1687,cstatus_csv_dumper_1687);
    fifo_csv_dumper_1688 = new("./depth1688.csv");
    cstatus_csv_dumper_1688 = new("./chan_status1688.csv");
    fifo_monitor_1688 = new(fifo_csv_dumper_1688,fifo_intf_1688,cstatus_csv_dumper_1688);
    fifo_csv_dumper_1689 = new("./depth1689.csv");
    cstatus_csv_dumper_1689 = new("./chan_status1689.csv");
    fifo_monitor_1689 = new(fifo_csv_dumper_1689,fifo_intf_1689,cstatus_csv_dumper_1689);
    fifo_csv_dumper_1690 = new("./depth1690.csv");
    cstatus_csv_dumper_1690 = new("./chan_status1690.csv");
    fifo_monitor_1690 = new(fifo_csv_dumper_1690,fifo_intf_1690,cstatus_csv_dumper_1690);
    fifo_csv_dumper_1691 = new("./depth1691.csv");
    cstatus_csv_dumper_1691 = new("./chan_status1691.csv");
    fifo_monitor_1691 = new(fifo_csv_dumper_1691,fifo_intf_1691,cstatus_csv_dumper_1691);
    fifo_csv_dumper_1692 = new("./depth1692.csv");
    cstatus_csv_dumper_1692 = new("./chan_status1692.csv");
    fifo_monitor_1692 = new(fifo_csv_dumper_1692,fifo_intf_1692,cstatus_csv_dumper_1692);
    fifo_csv_dumper_1693 = new("./depth1693.csv");
    cstatus_csv_dumper_1693 = new("./chan_status1693.csv");
    fifo_monitor_1693 = new(fifo_csv_dumper_1693,fifo_intf_1693,cstatus_csv_dumper_1693);
    fifo_csv_dumper_1694 = new("./depth1694.csv");
    cstatus_csv_dumper_1694 = new("./chan_status1694.csv");
    fifo_monitor_1694 = new(fifo_csv_dumper_1694,fifo_intf_1694,cstatus_csv_dumper_1694);
    fifo_csv_dumper_1695 = new("./depth1695.csv");
    cstatus_csv_dumper_1695 = new("./chan_status1695.csv");
    fifo_monitor_1695 = new(fifo_csv_dumper_1695,fifo_intf_1695,cstatus_csv_dumper_1695);
    fifo_csv_dumper_1696 = new("./depth1696.csv");
    cstatus_csv_dumper_1696 = new("./chan_status1696.csv");
    fifo_monitor_1696 = new(fifo_csv_dumper_1696,fifo_intf_1696,cstatus_csv_dumper_1696);
    fifo_csv_dumper_1697 = new("./depth1697.csv");
    cstatus_csv_dumper_1697 = new("./chan_status1697.csv");
    fifo_monitor_1697 = new(fifo_csv_dumper_1697,fifo_intf_1697,cstatus_csv_dumper_1697);
    fifo_csv_dumper_1698 = new("./depth1698.csv");
    cstatus_csv_dumper_1698 = new("./chan_status1698.csv");
    fifo_monitor_1698 = new(fifo_csv_dumper_1698,fifo_intf_1698,cstatus_csv_dumper_1698);
    fifo_csv_dumper_1699 = new("./depth1699.csv");
    cstatus_csv_dumper_1699 = new("./chan_status1699.csv");
    fifo_monitor_1699 = new(fifo_csv_dumper_1699,fifo_intf_1699,cstatus_csv_dumper_1699);
    fifo_csv_dumper_1700 = new("./depth1700.csv");
    cstatus_csv_dumper_1700 = new("./chan_status1700.csv");
    fifo_monitor_1700 = new(fifo_csv_dumper_1700,fifo_intf_1700,cstatus_csv_dumper_1700);
    fifo_csv_dumper_1701 = new("./depth1701.csv");
    cstatus_csv_dumper_1701 = new("./chan_status1701.csv");
    fifo_monitor_1701 = new(fifo_csv_dumper_1701,fifo_intf_1701,cstatus_csv_dumper_1701);
    fifo_csv_dumper_1702 = new("./depth1702.csv");
    cstatus_csv_dumper_1702 = new("./chan_status1702.csv");
    fifo_monitor_1702 = new(fifo_csv_dumper_1702,fifo_intf_1702,cstatus_csv_dumper_1702);
    fifo_csv_dumper_1703 = new("./depth1703.csv");
    cstatus_csv_dumper_1703 = new("./chan_status1703.csv");
    fifo_monitor_1703 = new(fifo_csv_dumper_1703,fifo_intf_1703,cstatus_csv_dumper_1703);
    fifo_csv_dumper_1704 = new("./depth1704.csv");
    cstatus_csv_dumper_1704 = new("./chan_status1704.csv");
    fifo_monitor_1704 = new(fifo_csv_dumper_1704,fifo_intf_1704,cstatus_csv_dumper_1704);
    fifo_csv_dumper_1705 = new("./depth1705.csv");
    cstatus_csv_dumper_1705 = new("./chan_status1705.csv");
    fifo_monitor_1705 = new(fifo_csv_dumper_1705,fifo_intf_1705,cstatus_csv_dumper_1705);
    fifo_csv_dumper_1706 = new("./depth1706.csv");
    cstatus_csv_dumper_1706 = new("./chan_status1706.csv");
    fifo_monitor_1706 = new(fifo_csv_dumper_1706,fifo_intf_1706,cstatus_csv_dumper_1706);
    fifo_csv_dumper_1707 = new("./depth1707.csv");
    cstatus_csv_dumper_1707 = new("./chan_status1707.csv");
    fifo_monitor_1707 = new(fifo_csv_dumper_1707,fifo_intf_1707,cstatus_csv_dumper_1707);
    fifo_csv_dumper_1708 = new("./depth1708.csv");
    cstatus_csv_dumper_1708 = new("./chan_status1708.csv");
    fifo_monitor_1708 = new(fifo_csv_dumper_1708,fifo_intf_1708,cstatus_csv_dumper_1708);
    fifo_csv_dumper_1709 = new("./depth1709.csv");
    cstatus_csv_dumper_1709 = new("./chan_status1709.csv");
    fifo_monitor_1709 = new(fifo_csv_dumper_1709,fifo_intf_1709,cstatus_csv_dumper_1709);
    fifo_csv_dumper_1710 = new("./depth1710.csv");
    cstatus_csv_dumper_1710 = new("./chan_status1710.csv");
    fifo_monitor_1710 = new(fifo_csv_dumper_1710,fifo_intf_1710,cstatus_csv_dumper_1710);
    fifo_csv_dumper_1711 = new("./depth1711.csv");
    cstatus_csv_dumper_1711 = new("./chan_status1711.csv");
    fifo_monitor_1711 = new(fifo_csv_dumper_1711,fifo_intf_1711,cstatus_csv_dumper_1711);
    fifo_csv_dumper_1712 = new("./depth1712.csv");
    cstatus_csv_dumper_1712 = new("./chan_status1712.csv");
    fifo_monitor_1712 = new(fifo_csv_dumper_1712,fifo_intf_1712,cstatus_csv_dumper_1712);
    fifo_csv_dumper_1713 = new("./depth1713.csv");
    cstatus_csv_dumper_1713 = new("./chan_status1713.csv");
    fifo_monitor_1713 = new(fifo_csv_dumper_1713,fifo_intf_1713,cstatus_csv_dumper_1713);
    fifo_csv_dumper_1714 = new("./depth1714.csv");
    cstatus_csv_dumper_1714 = new("./chan_status1714.csv");
    fifo_monitor_1714 = new(fifo_csv_dumper_1714,fifo_intf_1714,cstatus_csv_dumper_1714);
    fifo_csv_dumper_1715 = new("./depth1715.csv");
    cstatus_csv_dumper_1715 = new("./chan_status1715.csv");
    fifo_monitor_1715 = new(fifo_csv_dumper_1715,fifo_intf_1715,cstatus_csv_dumper_1715);
    fifo_csv_dumper_1716 = new("./depth1716.csv");
    cstatus_csv_dumper_1716 = new("./chan_status1716.csv");
    fifo_monitor_1716 = new(fifo_csv_dumper_1716,fifo_intf_1716,cstatus_csv_dumper_1716);
    fifo_csv_dumper_1717 = new("./depth1717.csv");
    cstatus_csv_dumper_1717 = new("./chan_status1717.csv");
    fifo_monitor_1717 = new(fifo_csv_dumper_1717,fifo_intf_1717,cstatus_csv_dumper_1717);
    fifo_csv_dumper_1718 = new("./depth1718.csv");
    cstatus_csv_dumper_1718 = new("./chan_status1718.csv");
    fifo_monitor_1718 = new(fifo_csv_dumper_1718,fifo_intf_1718,cstatus_csv_dumper_1718);
    fifo_csv_dumper_1719 = new("./depth1719.csv");
    cstatus_csv_dumper_1719 = new("./chan_status1719.csv");
    fifo_monitor_1719 = new(fifo_csv_dumper_1719,fifo_intf_1719,cstatus_csv_dumper_1719);
    fifo_csv_dumper_1720 = new("./depth1720.csv");
    cstatus_csv_dumper_1720 = new("./chan_status1720.csv");
    fifo_monitor_1720 = new(fifo_csv_dumper_1720,fifo_intf_1720,cstatus_csv_dumper_1720);
    fifo_csv_dumper_1721 = new("./depth1721.csv");
    cstatus_csv_dumper_1721 = new("./chan_status1721.csv");
    fifo_monitor_1721 = new(fifo_csv_dumper_1721,fifo_intf_1721,cstatus_csv_dumper_1721);
    fifo_csv_dumper_1722 = new("./depth1722.csv");
    cstatus_csv_dumper_1722 = new("./chan_status1722.csv");
    fifo_monitor_1722 = new(fifo_csv_dumper_1722,fifo_intf_1722,cstatus_csv_dumper_1722);
    fifo_csv_dumper_1723 = new("./depth1723.csv");
    cstatus_csv_dumper_1723 = new("./chan_status1723.csv");
    fifo_monitor_1723 = new(fifo_csv_dumper_1723,fifo_intf_1723,cstatus_csv_dumper_1723);
    fifo_csv_dumper_1724 = new("./depth1724.csv");
    cstatus_csv_dumper_1724 = new("./chan_status1724.csv");
    fifo_monitor_1724 = new(fifo_csv_dumper_1724,fifo_intf_1724,cstatus_csv_dumper_1724);
    fifo_csv_dumper_1725 = new("./depth1725.csv");
    cstatus_csv_dumper_1725 = new("./chan_status1725.csv");
    fifo_monitor_1725 = new(fifo_csv_dumper_1725,fifo_intf_1725,cstatus_csv_dumper_1725);
    fifo_csv_dumper_1726 = new("./depth1726.csv");
    cstatus_csv_dumper_1726 = new("./chan_status1726.csv");
    fifo_monitor_1726 = new(fifo_csv_dumper_1726,fifo_intf_1726,cstatus_csv_dumper_1726);
    fifo_csv_dumper_1727 = new("./depth1727.csv");
    cstatus_csv_dumper_1727 = new("./chan_status1727.csv");
    fifo_monitor_1727 = new(fifo_csv_dumper_1727,fifo_intf_1727,cstatus_csv_dumper_1727);
    fifo_csv_dumper_1728 = new("./depth1728.csv");
    cstatus_csv_dumper_1728 = new("./chan_status1728.csv");
    fifo_monitor_1728 = new(fifo_csv_dumper_1728,fifo_intf_1728,cstatus_csv_dumper_1728);
    fifo_csv_dumper_1729 = new("./depth1729.csv");
    cstatus_csv_dumper_1729 = new("./chan_status1729.csv");
    fifo_monitor_1729 = new(fifo_csv_dumper_1729,fifo_intf_1729,cstatus_csv_dumper_1729);
    fifo_csv_dumper_1730 = new("./depth1730.csv");
    cstatus_csv_dumper_1730 = new("./chan_status1730.csv");
    fifo_monitor_1730 = new(fifo_csv_dumper_1730,fifo_intf_1730,cstatus_csv_dumper_1730);
    fifo_csv_dumper_1731 = new("./depth1731.csv");
    cstatus_csv_dumper_1731 = new("./chan_status1731.csv");
    fifo_monitor_1731 = new(fifo_csv_dumper_1731,fifo_intf_1731,cstatus_csv_dumper_1731);
    fifo_csv_dumper_1732 = new("./depth1732.csv");
    cstatus_csv_dumper_1732 = new("./chan_status1732.csv");
    fifo_monitor_1732 = new(fifo_csv_dumper_1732,fifo_intf_1732,cstatus_csv_dumper_1732);
    fifo_csv_dumper_1733 = new("./depth1733.csv");
    cstatus_csv_dumper_1733 = new("./chan_status1733.csv");
    fifo_monitor_1733 = new(fifo_csv_dumper_1733,fifo_intf_1733,cstatus_csv_dumper_1733);
    fifo_csv_dumper_1734 = new("./depth1734.csv");
    cstatus_csv_dumper_1734 = new("./chan_status1734.csv");
    fifo_monitor_1734 = new(fifo_csv_dumper_1734,fifo_intf_1734,cstatus_csv_dumper_1734);
    fifo_csv_dumper_1735 = new("./depth1735.csv");
    cstatus_csv_dumper_1735 = new("./chan_status1735.csv");
    fifo_monitor_1735 = new(fifo_csv_dumper_1735,fifo_intf_1735,cstatus_csv_dumper_1735);
    fifo_csv_dumper_1736 = new("./depth1736.csv");
    cstatus_csv_dumper_1736 = new("./chan_status1736.csv");
    fifo_monitor_1736 = new(fifo_csv_dumper_1736,fifo_intf_1736,cstatus_csv_dumper_1736);
    fifo_csv_dumper_1737 = new("./depth1737.csv");
    cstatus_csv_dumper_1737 = new("./chan_status1737.csv");
    fifo_monitor_1737 = new(fifo_csv_dumper_1737,fifo_intf_1737,cstatus_csv_dumper_1737);
    fifo_csv_dumper_1738 = new("./depth1738.csv");
    cstatus_csv_dumper_1738 = new("./chan_status1738.csv");
    fifo_monitor_1738 = new(fifo_csv_dumper_1738,fifo_intf_1738,cstatus_csv_dumper_1738);
    fifo_csv_dumper_1739 = new("./depth1739.csv");
    cstatus_csv_dumper_1739 = new("./chan_status1739.csv");
    fifo_monitor_1739 = new(fifo_csv_dumper_1739,fifo_intf_1739,cstatus_csv_dumper_1739);
    fifo_csv_dumper_1740 = new("./depth1740.csv");
    cstatus_csv_dumper_1740 = new("./chan_status1740.csv");
    fifo_monitor_1740 = new(fifo_csv_dumper_1740,fifo_intf_1740,cstatus_csv_dumper_1740);
    fifo_csv_dumper_1741 = new("./depth1741.csv");
    cstatus_csv_dumper_1741 = new("./chan_status1741.csv");
    fifo_monitor_1741 = new(fifo_csv_dumper_1741,fifo_intf_1741,cstatus_csv_dumper_1741);
    fifo_csv_dumper_1742 = new("./depth1742.csv");
    cstatus_csv_dumper_1742 = new("./chan_status1742.csv");
    fifo_monitor_1742 = new(fifo_csv_dumper_1742,fifo_intf_1742,cstatus_csv_dumper_1742);
    fifo_csv_dumper_1743 = new("./depth1743.csv");
    cstatus_csv_dumper_1743 = new("./chan_status1743.csv");
    fifo_monitor_1743 = new(fifo_csv_dumper_1743,fifo_intf_1743,cstatus_csv_dumper_1743);
    fifo_csv_dumper_1744 = new("./depth1744.csv");
    cstatus_csv_dumper_1744 = new("./chan_status1744.csv");
    fifo_monitor_1744 = new(fifo_csv_dumper_1744,fifo_intf_1744,cstatus_csv_dumper_1744);
    fifo_csv_dumper_1745 = new("./depth1745.csv");
    cstatus_csv_dumper_1745 = new("./chan_status1745.csv");
    fifo_monitor_1745 = new(fifo_csv_dumper_1745,fifo_intf_1745,cstatus_csv_dumper_1745);
    fifo_csv_dumper_1746 = new("./depth1746.csv");
    cstatus_csv_dumper_1746 = new("./chan_status1746.csv");
    fifo_monitor_1746 = new(fifo_csv_dumper_1746,fifo_intf_1746,cstatus_csv_dumper_1746);
    fifo_csv_dumper_1747 = new("./depth1747.csv");
    cstatus_csv_dumper_1747 = new("./chan_status1747.csv");
    fifo_monitor_1747 = new(fifo_csv_dumper_1747,fifo_intf_1747,cstatus_csv_dumper_1747);
    fifo_csv_dumper_1748 = new("./depth1748.csv");
    cstatus_csv_dumper_1748 = new("./chan_status1748.csv");
    fifo_monitor_1748 = new(fifo_csv_dumper_1748,fifo_intf_1748,cstatus_csv_dumper_1748);
    fifo_csv_dumper_1749 = new("./depth1749.csv");
    cstatus_csv_dumper_1749 = new("./chan_status1749.csv");
    fifo_monitor_1749 = new(fifo_csv_dumper_1749,fifo_intf_1749,cstatus_csv_dumper_1749);
    fifo_csv_dumper_1750 = new("./depth1750.csv");
    cstatus_csv_dumper_1750 = new("./chan_status1750.csv");
    fifo_monitor_1750 = new(fifo_csv_dumper_1750,fifo_intf_1750,cstatus_csv_dumper_1750);
    fifo_csv_dumper_1751 = new("./depth1751.csv");
    cstatus_csv_dumper_1751 = new("./chan_status1751.csv");
    fifo_monitor_1751 = new(fifo_csv_dumper_1751,fifo_intf_1751,cstatus_csv_dumper_1751);
    fifo_csv_dumper_1752 = new("./depth1752.csv");
    cstatus_csv_dumper_1752 = new("./chan_status1752.csv");
    fifo_monitor_1752 = new(fifo_csv_dumper_1752,fifo_intf_1752,cstatus_csv_dumper_1752);
    fifo_csv_dumper_1753 = new("./depth1753.csv");
    cstatus_csv_dumper_1753 = new("./chan_status1753.csv");
    fifo_monitor_1753 = new(fifo_csv_dumper_1753,fifo_intf_1753,cstatus_csv_dumper_1753);
    fifo_csv_dumper_1754 = new("./depth1754.csv");
    cstatus_csv_dumper_1754 = new("./chan_status1754.csv");
    fifo_monitor_1754 = new(fifo_csv_dumper_1754,fifo_intf_1754,cstatus_csv_dumper_1754);
    fifo_csv_dumper_1755 = new("./depth1755.csv");
    cstatus_csv_dumper_1755 = new("./chan_status1755.csv");
    fifo_monitor_1755 = new(fifo_csv_dumper_1755,fifo_intf_1755,cstatus_csv_dumper_1755);
    fifo_csv_dumper_1756 = new("./depth1756.csv");
    cstatus_csv_dumper_1756 = new("./chan_status1756.csv");
    fifo_monitor_1756 = new(fifo_csv_dumper_1756,fifo_intf_1756,cstatus_csv_dumper_1756);
    fifo_csv_dumper_1757 = new("./depth1757.csv");
    cstatus_csv_dumper_1757 = new("./chan_status1757.csv");
    fifo_monitor_1757 = new(fifo_csv_dumper_1757,fifo_intf_1757,cstatus_csv_dumper_1757);
    fifo_csv_dumper_1758 = new("./depth1758.csv");
    cstatus_csv_dumper_1758 = new("./chan_status1758.csv");
    fifo_monitor_1758 = new(fifo_csv_dumper_1758,fifo_intf_1758,cstatus_csv_dumper_1758);
    fifo_csv_dumper_1759 = new("./depth1759.csv");
    cstatus_csv_dumper_1759 = new("./chan_status1759.csv");
    fifo_monitor_1759 = new(fifo_csv_dumper_1759,fifo_intf_1759,cstatus_csv_dumper_1759);
    fifo_csv_dumper_1760 = new("./depth1760.csv");
    cstatus_csv_dumper_1760 = new("./chan_status1760.csv");
    fifo_monitor_1760 = new(fifo_csv_dumper_1760,fifo_intf_1760,cstatus_csv_dumper_1760);
    fifo_csv_dumper_1761 = new("./depth1761.csv");
    cstatus_csv_dumper_1761 = new("./chan_status1761.csv");
    fifo_monitor_1761 = new(fifo_csv_dumper_1761,fifo_intf_1761,cstatus_csv_dumper_1761);
    fifo_csv_dumper_1762 = new("./depth1762.csv");
    cstatus_csv_dumper_1762 = new("./chan_status1762.csv");
    fifo_monitor_1762 = new(fifo_csv_dumper_1762,fifo_intf_1762,cstatus_csv_dumper_1762);
    fifo_csv_dumper_1763 = new("./depth1763.csv");
    cstatus_csv_dumper_1763 = new("./chan_status1763.csv");
    fifo_monitor_1763 = new(fifo_csv_dumper_1763,fifo_intf_1763,cstatus_csv_dumper_1763);
    fifo_csv_dumper_1764 = new("./depth1764.csv");
    cstatus_csv_dumper_1764 = new("./chan_status1764.csv");
    fifo_monitor_1764 = new(fifo_csv_dumper_1764,fifo_intf_1764,cstatus_csv_dumper_1764);
    fifo_csv_dumper_1765 = new("./depth1765.csv");
    cstatus_csv_dumper_1765 = new("./chan_status1765.csv");
    fifo_monitor_1765 = new(fifo_csv_dumper_1765,fifo_intf_1765,cstatus_csv_dumper_1765);
    fifo_csv_dumper_1766 = new("./depth1766.csv");
    cstatus_csv_dumper_1766 = new("./chan_status1766.csv");
    fifo_monitor_1766 = new(fifo_csv_dumper_1766,fifo_intf_1766,cstatus_csv_dumper_1766);
    fifo_csv_dumper_1767 = new("./depth1767.csv");
    cstatus_csv_dumper_1767 = new("./chan_status1767.csv");
    fifo_monitor_1767 = new(fifo_csv_dumper_1767,fifo_intf_1767,cstatus_csv_dumper_1767);
    fifo_csv_dumper_1768 = new("./depth1768.csv");
    cstatus_csv_dumper_1768 = new("./chan_status1768.csv");
    fifo_monitor_1768 = new(fifo_csv_dumper_1768,fifo_intf_1768,cstatus_csv_dumper_1768);
    fifo_csv_dumper_1769 = new("./depth1769.csv");
    cstatus_csv_dumper_1769 = new("./chan_status1769.csv");
    fifo_monitor_1769 = new(fifo_csv_dumper_1769,fifo_intf_1769,cstatus_csv_dumper_1769);
    fifo_csv_dumper_1770 = new("./depth1770.csv");
    cstatus_csv_dumper_1770 = new("./chan_status1770.csv");
    fifo_monitor_1770 = new(fifo_csv_dumper_1770,fifo_intf_1770,cstatus_csv_dumper_1770);
    fifo_csv_dumper_1771 = new("./depth1771.csv");
    cstatus_csv_dumper_1771 = new("./chan_status1771.csv");
    fifo_monitor_1771 = new(fifo_csv_dumper_1771,fifo_intf_1771,cstatus_csv_dumper_1771);
    fifo_csv_dumper_1772 = new("./depth1772.csv");
    cstatus_csv_dumper_1772 = new("./chan_status1772.csv");
    fifo_monitor_1772 = new(fifo_csv_dumper_1772,fifo_intf_1772,cstatus_csv_dumper_1772);
    fifo_csv_dumper_1773 = new("./depth1773.csv");
    cstatus_csv_dumper_1773 = new("./chan_status1773.csv");
    fifo_monitor_1773 = new(fifo_csv_dumper_1773,fifo_intf_1773,cstatus_csv_dumper_1773);
    fifo_csv_dumper_1774 = new("./depth1774.csv");
    cstatus_csv_dumper_1774 = new("./chan_status1774.csv");
    fifo_monitor_1774 = new(fifo_csv_dumper_1774,fifo_intf_1774,cstatus_csv_dumper_1774);
    fifo_csv_dumper_1775 = new("./depth1775.csv");
    cstatus_csv_dumper_1775 = new("./chan_status1775.csv");
    fifo_monitor_1775 = new(fifo_csv_dumper_1775,fifo_intf_1775,cstatus_csv_dumper_1775);
    fifo_csv_dumper_1776 = new("./depth1776.csv");
    cstatus_csv_dumper_1776 = new("./chan_status1776.csv");
    fifo_monitor_1776 = new(fifo_csv_dumper_1776,fifo_intf_1776,cstatus_csv_dumper_1776);
    fifo_csv_dumper_1777 = new("./depth1777.csv");
    cstatus_csv_dumper_1777 = new("./chan_status1777.csv");
    fifo_monitor_1777 = new(fifo_csv_dumper_1777,fifo_intf_1777,cstatus_csv_dumper_1777);
    fifo_csv_dumper_1778 = new("./depth1778.csv");
    cstatus_csv_dumper_1778 = new("./chan_status1778.csv");
    fifo_monitor_1778 = new(fifo_csv_dumper_1778,fifo_intf_1778,cstatus_csv_dumper_1778);
    fifo_csv_dumper_1779 = new("./depth1779.csv");
    cstatus_csv_dumper_1779 = new("./chan_status1779.csv");
    fifo_monitor_1779 = new(fifo_csv_dumper_1779,fifo_intf_1779,cstatus_csv_dumper_1779);
    fifo_csv_dumper_1780 = new("./depth1780.csv");
    cstatus_csv_dumper_1780 = new("./chan_status1780.csv");
    fifo_monitor_1780 = new(fifo_csv_dumper_1780,fifo_intf_1780,cstatus_csv_dumper_1780);
    fifo_csv_dumper_1781 = new("./depth1781.csv");
    cstatus_csv_dumper_1781 = new("./chan_status1781.csv");
    fifo_monitor_1781 = new(fifo_csv_dumper_1781,fifo_intf_1781,cstatus_csv_dumper_1781);
    fifo_csv_dumper_1782 = new("./depth1782.csv");
    cstatus_csv_dumper_1782 = new("./chan_status1782.csv");
    fifo_monitor_1782 = new(fifo_csv_dumper_1782,fifo_intf_1782,cstatus_csv_dumper_1782);
    fifo_csv_dumper_1783 = new("./depth1783.csv");
    cstatus_csv_dumper_1783 = new("./chan_status1783.csv");
    fifo_monitor_1783 = new(fifo_csv_dumper_1783,fifo_intf_1783,cstatus_csv_dumper_1783);
    fifo_csv_dumper_1784 = new("./depth1784.csv");
    cstatus_csv_dumper_1784 = new("./chan_status1784.csv");
    fifo_monitor_1784 = new(fifo_csv_dumper_1784,fifo_intf_1784,cstatus_csv_dumper_1784);
    fifo_csv_dumper_1785 = new("./depth1785.csv");
    cstatus_csv_dumper_1785 = new("./chan_status1785.csv");
    fifo_monitor_1785 = new(fifo_csv_dumper_1785,fifo_intf_1785,cstatus_csv_dumper_1785);
    fifo_csv_dumper_1786 = new("./depth1786.csv");
    cstatus_csv_dumper_1786 = new("./chan_status1786.csv");
    fifo_monitor_1786 = new(fifo_csv_dumper_1786,fifo_intf_1786,cstatus_csv_dumper_1786);
    fifo_csv_dumper_1787 = new("./depth1787.csv");
    cstatus_csv_dumper_1787 = new("./chan_status1787.csv");
    fifo_monitor_1787 = new(fifo_csv_dumper_1787,fifo_intf_1787,cstatus_csv_dumper_1787);
    fifo_csv_dumper_1788 = new("./depth1788.csv");
    cstatus_csv_dumper_1788 = new("./chan_status1788.csv");
    fifo_monitor_1788 = new(fifo_csv_dumper_1788,fifo_intf_1788,cstatus_csv_dumper_1788);
    fifo_csv_dumper_1789 = new("./depth1789.csv");
    cstatus_csv_dumper_1789 = new("./chan_status1789.csv");
    fifo_monitor_1789 = new(fifo_csv_dumper_1789,fifo_intf_1789,cstatus_csv_dumper_1789);
    fifo_csv_dumper_1790 = new("./depth1790.csv");
    cstatus_csv_dumper_1790 = new("./chan_status1790.csv");
    fifo_monitor_1790 = new(fifo_csv_dumper_1790,fifo_intf_1790,cstatus_csv_dumper_1790);
    fifo_csv_dumper_1791 = new("./depth1791.csv");
    cstatus_csv_dumper_1791 = new("./chan_status1791.csv");
    fifo_monitor_1791 = new(fifo_csv_dumper_1791,fifo_intf_1791,cstatus_csv_dumper_1791);
    fifo_csv_dumper_1792 = new("./depth1792.csv");
    cstatus_csv_dumper_1792 = new("./chan_status1792.csv");
    fifo_monitor_1792 = new(fifo_csv_dumper_1792,fifo_intf_1792,cstatus_csv_dumper_1792);
    fifo_csv_dumper_1793 = new("./depth1793.csv");
    cstatus_csv_dumper_1793 = new("./chan_status1793.csv");
    fifo_monitor_1793 = new(fifo_csv_dumper_1793,fifo_intf_1793,cstatus_csv_dumper_1793);
    fifo_csv_dumper_1794 = new("./depth1794.csv");
    cstatus_csv_dumper_1794 = new("./chan_status1794.csv");
    fifo_monitor_1794 = new(fifo_csv_dumper_1794,fifo_intf_1794,cstatus_csv_dumper_1794);
    fifo_csv_dumper_1795 = new("./depth1795.csv");
    cstatus_csv_dumper_1795 = new("./chan_status1795.csv");
    fifo_monitor_1795 = new(fifo_csv_dumper_1795,fifo_intf_1795,cstatus_csv_dumper_1795);
    fifo_csv_dumper_1796 = new("./depth1796.csv");
    cstatus_csv_dumper_1796 = new("./chan_status1796.csv");
    fifo_monitor_1796 = new(fifo_csv_dumper_1796,fifo_intf_1796,cstatus_csv_dumper_1796);
    fifo_csv_dumper_1797 = new("./depth1797.csv");
    cstatus_csv_dumper_1797 = new("./chan_status1797.csv");
    fifo_monitor_1797 = new(fifo_csv_dumper_1797,fifo_intf_1797,cstatus_csv_dumper_1797);
    fifo_csv_dumper_1798 = new("./depth1798.csv");
    cstatus_csv_dumper_1798 = new("./chan_status1798.csv");
    fifo_monitor_1798 = new(fifo_csv_dumper_1798,fifo_intf_1798,cstatus_csv_dumper_1798);
    fifo_csv_dumper_1799 = new("./depth1799.csv");
    cstatus_csv_dumper_1799 = new("./chan_status1799.csv");
    fifo_monitor_1799 = new(fifo_csv_dumper_1799,fifo_intf_1799,cstatus_csv_dumper_1799);
    fifo_csv_dumper_1800 = new("./depth1800.csv");
    cstatus_csv_dumper_1800 = new("./chan_status1800.csv");
    fifo_monitor_1800 = new(fifo_csv_dumper_1800,fifo_intf_1800,cstatus_csv_dumper_1800);
    fifo_csv_dumper_1801 = new("./depth1801.csv");
    cstatus_csv_dumper_1801 = new("./chan_status1801.csv");
    fifo_monitor_1801 = new(fifo_csv_dumper_1801,fifo_intf_1801,cstatus_csv_dumper_1801);
    fifo_csv_dumper_1802 = new("./depth1802.csv");
    cstatus_csv_dumper_1802 = new("./chan_status1802.csv");
    fifo_monitor_1802 = new(fifo_csv_dumper_1802,fifo_intf_1802,cstatus_csv_dumper_1802);
    fifo_csv_dumper_1803 = new("./depth1803.csv");
    cstatus_csv_dumper_1803 = new("./chan_status1803.csv");
    fifo_monitor_1803 = new(fifo_csv_dumper_1803,fifo_intf_1803,cstatus_csv_dumper_1803);
    fifo_csv_dumper_1804 = new("./depth1804.csv");
    cstatus_csv_dumper_1804 = new("./chan_status1804.csv");
    fifo_monitor_1804 = new(fifo_csv_dumper_1804,fifo_intf_1804,cstatus_csv_dumper_1804);
    fifo_csv_dumper_1805 = new("./depth1805.csv");
    cstatus_csv_dumper_1805 = new("./chan_status1805.csv");
    fifo_monitor_1805 = new(fifo_csv_dumper_1805,fifo_intf_1805,cstatus_csv_dumper_1805);
    fifo_csv_dumper_1806 = new("./depth1806.csv");
    cstatus_csv_dumper_1806 = new("./chan_status1806.csv");
    fifo_monitor_1806 = new(fifo_csv_dumper_1806,fifo_intf_1806,cstatus_csv_dumper_1806);
    fifo_csv_dumper_1807 = new("./depth1807.csv");
    cstatus_csv_dumper_1807 = new("./chan_status1807.csv");
    fifo_monitor_1807 = new(fifo_csv_dumper_1807,fifo_intf_1807,cstatus_csv_dumper_1807);
    fifo_csv_dumper_1808 = new("./depth1808.csv");
    cstatus_csv_dumper_1808 = new("./chan_status1808.csv");
    fifo_monitor_1808 = new(fifo_csv_dumper_1808,fifo_intf_1808,cstatus_csv_dumper_1808);
    fifo_csv_dumper_1809 = new("./depth1809.csv");
    cstatus_csv_dumper_1809 = new("./chan_status1809.csv");
    fifo_monitor_1809 = new(fifo_csv_dumper_1809,fifo_intf_1809,cstatus_csv_dumper_1809);
    fifo_csv_dumper_1810 = new("./depth1810.csv");
    cstatus_csv_dumper_1810 = new("./chan_status1810.csv");
    fifo_monitor_1810 = new(fifo_csv_dumper_1810,fifo_intf_1810,cstatus_csv_dumper_1810);
    fifo_csv_dumper_1811 = new("./depth1811.csv");
    cstatus_csv_dumper_1811 = new("./chan_status1811.csv");
    fifo_monitor_1811 = new(fifo_csv_dumper_1811,fifo_intf_1811,cstatus_csv_dumper_1811);
    fifo_csv_dumper_1812 = new("./depth1812.csv");
    cstatus_csv_dumper_1812 = new("./chan_status1812.csv");
    fifo_monitor_1812 = new(fifo_csv_dumper_1812,fifo_intf_1812,cstatus_csv_dumper_1812);
    fifo_csv_dumper_1813 = new("./depth1813.csv");
    cstatus_csv_dumper_1813 = new("./chan_status1813.csv");
    fifo_monitor_1813 = new(fifo_csv_dumper_1813,fifo_intf_1813,cstatus_csv_dumper_1813);
    fifo_csv_dumper_1814 = new("./depth1814.csv");
    cstatus_csv_dumper_1814 = new("./chan_status1814.csv");
    fifo_monitor_1814 = new(fifo_csv_dumper_1814,fifo_intf_1814,cstatus_csv_dumper_1814);
    fifo_csv_dumper_1815 = new("./depth1815.csv");
    cstatus_csv_dumper_1815 = new("./chan_status1815.csv");
    fifo_monitor_1815 = new(fifo_csv_dumper_1815,fifo_intf_1815,cstatus_csv_dumper_1815);
    fifo_csv_dumper_1816 = new("./depth1816.csv");
    cstatus_csv_dumper_1816 = new("./chan_status1816.csv");
    fifo_monitor_1816 = new(fifo_csv_dumper_1816,fifo_intf_1816,cstatus_csv_dumper_1816);
    fifo_csv_dumper_1817 = new("./depth1817.csv");
    cstatus_csv_dumper_1817 = new("./chan_status1817.csv");
    fifo_monitor_1817 = new(fifo_csv_dumper_1817,fifo_intf_1817,cstatus_csv_dumper_1817);
    fifo_csv_dumper_1818 = new("./depth1818.csv");
    cstatus_csv_dumper_1818 = new("./chan_status1818.csv");
    fifo_monitor_1818 = new(fifo_csv_dumper_1818,fifo_intf_1818,cstatus_csv_dumper_1818);
    fifo_csv_dumper_1819 = new("./depth1819.csv");
    cstatus_csv_dumper_1819 = new("./chan_status1819.csv");
    fifo_monitor_1819 = new(fifo_csv_dumper_1819,fifo_intf_1819,cstatus_csv_dumper_1819);
    fifo_csv_dumper_1820 = new("./depth1820.csv");
    cstatus_csv_dumper_1820 = new("./chan_status1820.csv");
    fifo_monitor_1820 = new(fifo_csv_dumper_1820,fifo_intf_1820,cstatus_csv_dumper_1820);
    fifo_csv_dumper_1821 = new("./depth1821.csv");
    cstatus_csv_dumper_1821 = new("./chan_status1821.csv");
    fifo_monitor_1821 = new(fifo_csv_dumper_1821,fifo_intf_1821,cstatus_csv_dumper_1821);
    fifo_csv_dumper_1822 = new("./depth1822.csv");
    cstatus_csv_dumper_1822 = new("./chan_status1822.csv");
    fifo_monitor_1822 = new(fifo_csv_dumper_1822,fifo_intf_1822,cstatus_csv_dumper_1822);
    fifo_csv_dumper_1823 = new("./depth1823.csv");
    cstatus_csv_dumper_1823 = new("./chan_status1823.csv");
    fifo_monitor_1823 = new(fifo_csv_dumper_1823,fifo_intf_1823,cstatus_csv_dumper_1823);
    fifo_csv_dumper_1824 = new("./depth1824.csv");
    cstatus_csv_dumper_1824 = new("./chan_status1824.csv");
    fifo_monitor_1824 = new(fifo_csv_dumper_1824,fifo_intf_1824,cstatus_csv_dumper_1824);
    fifo_csv_dumper_1825 = new("./depth1825.csv");
    cstatus_csv_dumper_1825 = new("./chan_status1825.csv");
    fifo_monitor_1825 = new(fifo_csv_dumper_1825,fifo_intf_1825,cstatus_csv_dumper_1825);
    fifo_csv_dumper_1826 = new("./depth1826.csv");
    cstatus_csv_dumper_1826 = new("./chan_status1826.csv");
    fifo_monitor_1826 = new(fifo_csv_dumper_1826,fifo_intf_1826,cstatus_csv_dumper_1826);
    fifo_csv_dumper_1827 = new("./depth1827.csv");
    cstatus_csv_dumper_1827 = new("./chan_status1827.csv");
    fifo_monitor_1827 = new(fifo_csv_dumper_1827,fifo_intf_1827,cstatus_csv_dumper_1827);
    fifo_csv_dumper_1828 = new("./depth1828.csv");
    cstatus_csv_dumper_1828 = new("./chan_status1828.csv");
    fifo_monitor_1828 = new(fifo_csv_dumper_1828,fifo_intf_1828,cstatus_csv_dumper_1828);
    fifo_csv_dumper_1829 = new("./depth1829.csv");
    cstatus_csv_dumper_1829 = new("./chan_status1829.csv");
    fifo_monitor_1829 = new(fifo_csv_dumper_1829,fifo_intf_1829,cstatus_csv_dumper_1829);
    fifo_csv_dumper_1830 = new("./depth1830.csv");
    cstatus_csv_dumper_1830 = new("./chan_status1830.csv");
    fifo_monitor_1830 = new(fifo_csv_dumper_1830,fifo_intf_1830,cstatus_csv_dumper_1830);
    fifo_csv_dumper_1831 = new("./depth1831.csv");
    cstatus_csv_dumper_1831 = new("./chan_status1831.csv");
    fifo_monitor_1831 = new(fifo_csv_dumper_1831,fifo_intf_1831,cstatus_csv_dumper_1831);
    fifo_csv_dumper_1832 = new("./depth1832.csv");
    cstatus_csv_dumper_1832 = new("./chan_status1832.csv");
    fifo_monitor_1832 = new(fifo_csv_dumper_1832,fifo_intf_1832,cstatus_csv_dumper_1832);
    fifo_csv_dumper_1833 = new("./depth1833.csv");
    cstatus_csv_dumper_1833 = new("./chan_status1833.csv");
    fifo_monitor_1833 = new(fifo_csv_dumper_1833,fifo_intf_1833,cstatus_csv_dumper_1833);
    fifo_csv_dumper_1834 = new("./depth1834.csv");
    cstatus_csv_dumper_1834 = new("./chan_status1834.csv");
    fifo_monitor_1834 = new(fifo_csv_dumper_1834,fifo_intf_1834,cstatus_csv_dumper_1834);
    fifo_csv_dumper_1835 = new("./depth1835.csv");
    cstatus_csv_dumper_1835 = new("./chan_status1835.csv");
    fifo_monitor_1835 = new(fifo_csv_dumper_1835,fifo_intf_1835,cstatus_csv_dumper_1835);
    fifo_csv_dumper_1836 = new("./depth1836.csv");
    cstatus_csv_dumper_1836 = new("./chan_status1836.csv");
    fifo_monitor_1836 = new(fifo_csv_dumper_1836,fifo_intf_1836,cstatus_csv_dumper_1836);
    fifo_csv_dumper_1837 = new("./depth1837.csv");
    cstatus_csv_dumper_1837 = new("./chan_status1837.csv");
    fifo_monitor_1837 = new(fifo_csv_dumper_1837,fifo_intf_1837,cstatus_csv_dumper_1837);
    fifo_csv_dumper_1838 = new("./depth1838.csv");
    cstatus_csv_dumper_1838 = new("./chan_status1838.csv");
    fifo_monitor_1838 = new(fifo_csv_dumper_1838,fifo_intf_1838,cstatus_csv_dumper_1838);
    fifo_csv_dumper_1839 = new("./depth1839.csv");
    cstatus_csv_dumper_1839 = new("./chan_status1839.csv");
    fifo_monitor_1839 = new(fifo_csv_dumper_1839,fifo_intf_1839,cstatus_csv_dumper_1839);
    fifo_csv_dumper_1840 = new("./depth1840.csv");
    cstatus_csv_dumper_1840 = new("./chan_status1840.csv");
    fifo_monitor_1840 = new(fifo_csv_dumper_1840,fifo_intf_1840,cstatus_csv_dumper_1840);
    fifo_csv_dumper_1841 = new("./depth1841.csv");
    cstatus_csv_dumper_1841 = new("./chan_status1841.csv");
    fifo_monitor_1841 = new(fifo_csv_dumper_1841,fifo_intf_1841,cstatus_csv_dumper_1841);
    fifo_csv_dumper_1842 = new("./depth1842.csv");
    cstatus_csv_dumper_1842 = new("./chan_status1842.csv");
    fifo_monitor_1842 = new(fifo_csv_dumper_1842,fifo_intf_1842,cstatus_csv_dumper_1842);
    fifo_csv_dumper_1843 = new("./depth1843.csv");
    cstatus_csv_dumper_1843 = new("./chan_status1843.csv");
    fifo_monitor_1843 = new(fifo_csv_dumper_1843,fifo_intf_1843,cstatus_csv_dumper_1843);
    fifo_csv_dumper_1844 = new("./depth1844.csv");
    cstatus_csv_dumper_1844 = new("./chan_status1844.csv");
    fifo_monitor_1844 = new(fifo_csv_dumper_1844,fifo_intf_1844,cstatus_csv_dumper_1844);
    fifo_csv_dumper_1845 = new("./depth1845.csv");
    cstatus_csv_dumper_1845 = new("./chan_status1845.csv");
    fifo_monitor_1845 = new(fifo_csv_dumper_1845,fifo_intf_1845,cstatus_csv_dumper_1845);
    fifo_csv_dumper_1846 = new("./depth1846.csv");
    cstatus_csv_dumper_1846 = new("./chan_status1846.csv");
    fifo_monitor_1846 = new(fifo_csv_dumper_1846,fifo_intf_1846,cstatus_csv_dumper_1846);
    fifo_csv_dumper_1847 = new("./depth1847.csv");
    cstatus_csv_dumper_1847 = new("./chan_status1847.csv");
    fifo_monitor_1847 = new(fifo_csv_dumper_1847,fifo_intf_1847,cstatus_csv_dumper_1847);
    fifo_csv_dumper_1848 = new("./depth1848.csv");
    cstatus_csv_dumper_1848 = new("./chan_status1848.csv");
    fifo_monitor_1848 = new(fifo_csv_dumper_1848,fifo_intf_1848,cstatus_csv_dumper_1848);
    fifo_csv_dumper_1849 = new("./depth1849.csv");
    cstatus_csv_dumper_1849 = new("./chan_status1849.csv");
    fifo_monitor_1849 = new(fifo_csv_dumper_1849,fifo_intf_1849,cstatus_csv_dumper_1849);
    fifo_csv_dumper_1850 = new("./depth1850.csv");
    cstatus_csv_dumper_1850 = new("./chan_status1850.csv");
    fifo_monitor_1850 = new(fifo_csv_dumper_1850,fifo_intf_1850,cstatus_csv_dumper_1850);
    fifo_csv_dumper_1851 = new("./depth1851.csv");
    cstatus_csv_dumper_1851 = new("./chan_status1851.csv");
    fifo_monitor_1851 = new(fifo_csv_dumper_1851,fifo_intf_1851,cstatus_csv_dumper_1851);
    fifo_csv_dumper_1852 = new("./depth1852.csv");
    cstatus_csv_dumper_1852 = new("./chan_status1852.csv");
    fifo_monitor_1852 = new(fifo_csv_dumper_1852,fifo_intf_1852,cstatus_csv_dumper_1852);
    fifo_csv_dumper_1853 = new("./depth1853.csv");
    cstatus_csv_dumper_1853 = new("./chan_status1853.csv");
    fifo_monitor_1853 = new(fifo_csv_dumper_1853,fifo_intf_1853,cstatus_csv_dumper_1853);
    fifo_csv_dumper_1854 = new("./depth1854.csv");
    cstatus_csv_dumper_1854 = new("./chan_status1854.csv");
    fifo_monitor_1854 = new(fifo_csv_dumper_1854,fifo_intf_1854,cstatus_csv_dumper_1854);
    fifo_csv_dumper_1855 = new("./depth1855.csv");
    cstatus_csv_dumper_1855 = new("./chan_status1855.csv");
    fifo_monitor_1855 = new(fifo_csv_dumper_1855,fifo_intf_1855,cstatus_csv_dumper_1855);
    fifo_csv_dumper_1856 = new("./depth1856.csv");
    cstatus_csv_dumper_1856 = new("./chan_status1856.csv");
    fifo_monitor_1856 = new(fifo_csv_dumper_1856,fifo_intf_1856,cstatus_csv_dumper_1856);
    fifo_csv_dumper_1857 = new("./depth1857.csv");
    cstatus_csv_dumper_1857 = new("./chan_status1857.csv");
    fifo_monitor_1857 = new(fifo_csv_dumper_1857,fifo_intf_1857,cstatus_csv_dumper_1857);
    fifo_csv_dumper_1858 = new("./depth1858.csv");
    cstatus_csv_dumper_1858 = new("./chan_status1858.csv");
    fifo_monitor_1858 = new(fifo_csv_dumper_1858,fifo_intf_1858,cstatus_csv_dumper_1858);
    fifo_csv_dumper_1859 = new("./depth1859.csv");
    cstatus_csv_dumper_1859 = new("./chan_status1859.csv");
    fifo_monitor_1859 = new(fifo_csv_dumper_1859,fifo_intf_1859,cstatus_csv_dumper_1859);
    fifo_csv_dumper_1860 = new("./depth1860.csv");
    cstatus_csv_dumper_1860 = new("./chan_status1860.csv");
    fifo_monitor_1860 = new(fifo_csv_dumper_1860,fifo_intf_1860,cstatus_csv_dumper_1860);
    fifo_csv_dumper_1861 = new("./depth1861.csv");
    cstatus_csv_dumper_1861 = new("./chan_status1861.csv");
    fifo_monitor_1861 = new(fifo_csv_dumper_1861,fifo_intf_1861,cstatus_csv_dumper_1861);
    fifo_csv_dumper_1862 = new("./depth1862.csv");
    cstatus_csv_dumper_1862 = new("./chan_status1862.csv");
    fifo_monitor_1862 = new(fifo_csv_dumper_1862,fifo_intf_1862,cstatus_csv_dumper_1862);
    fifo_csv_dumper_1863 = new("./depth1863.csv");
    cstatus_csv_dumper_1863 = new("./chan_status1863.csv");
    fifo_monitor_1863 = new(fifo_csv_dumper_1863,fifo_intf_1863,cstatus_csv_dumper_1863);
    fifo_csv_dumper_1864 = new("./depth1864.csv");
    cstatus_csv_dumper_1864 = new("./chan_status1864.csv");
    fifo_monitor_1864 = new(fifo_csv_dumper_1864,fifo_intf_1864,cstatus_csv_dumper_1864);
    fifo_csv_dumper_1865 = new("./depth1865.csv");
    cstatus_csv_dumper_1865 = new("./chan_status1865.csv");
    fifo_monitor_1865 = new(fifo_csv_dumper_1865,fifo_intf_1865,cstatus_csv_dumper_1865);
    fifo_csv_dumper_1866 = new("./depth1866.csv");
    cstatus_csv_dumper_1866 = new("./chan_status1866.csv");
    fifo_monitor_1866 = new(fifo_csv_dumper_1866,fifo_intf_1866,cstatus_csv_dumper_1866);
    fifo_csv_dumper_1867 = new("./depth1867.csv");
    cstatus_csv_dumper_1867 = new("./chan_status1867.csv");
    fifo_monitor_1867 = new(fifo_csv_dumper_1867,fifo_intf_1867,cstatus_csv_dumper_1867);
    fifo_csv_dumper_1868 = new("./depth1868.csv");
    cstatus_csv_dumper_1868 = new("./chan_status1868.csv");
    fifo_monitor_1868 = new(fifo_csv_dumper_1868,fifo_intf_1868,cstatus_csv_dumper_1868);
    fifo_csv_dumper_1869 = new("./depth1869.csv");
    cstatus_csv_dumper_1869 = new("./chan_status1869.csv");
    fifo_monitor_1869 = new(fifo_csv_dumper_1869,fifo_intf_1869,cstatus_csv_dumper_1869);
    fifo_csv_dumper_1870 = new("./depth1870.csv");
    cstatus_csv_dumper_1870 = new("./chan_status1870.csv");
    fifo_monitor_1870 = new(fifo_csv_dumper_1870,fifo_intf_1870,cstatus_csv_dumper_1870);
    fifo_csv_dumper_1871 = new("./depth1871.csv");
    cstatus_csv_dumper_1871 = new("./chan_status1871.csv");
    fifo_monitor_1871 = new(fifo_csv_dumper_1871,fifo_intf_1871,cstatus_csv_dumper_1871);
    fifo_csv_dumper_1872 = new("./depth1872.csv");
    cstatus_csv_dumper_1872 = new("./chan_status1872.csv");
    fifo_monitor_1872 = new(fifo_csv_dumper_1872,fifo_intf_1872,cstatus_csv_dumper_1872);
    fifo_csv_dumper_1873 = new("./depth1873.csv");
    cstatus_csv_dumper_1873 = new("./chan_status1873.csv");
    fifo_monitor_1873 = new(fifo_csv_dumper_1873,fifo_intf_1873,cstatus_csv_dumper_1873);
    fifo_csv_dumper_1874 = new("./depth1874.csv");
    cstatus_csv_dumper_1874 = new("./chan_status1874.csv");
    fifo_monitor_1874 = new(fifo_csv_dumper_1874,fifo_intf_1874,cstatus_csv_dumper_1874);
    fifo_csv_dumper_1875 = new("./depth1875.csv");
    cstatus_csv_dumper_1875 = new("./chan_status1875.csv");
    fifo_monitor_1875 = new(fifo_csv_dumper_1875,fifo_intf_1875,cstatus_csv_dumper_1875);
    fifo_csv_dumper_1876 = new("./depth1876.csv");
    cstatus_csv_dumper_1876 = new("./chan_status1876.csv");
    fifo_monitor_1876 = new(fifo_csv_dumper_1876,fifo_intf_1876,cstatus_csv_dumper_1876);
    fifo_csv_dumper_1877 = new("./depth1877.csv");
    cstatus_csv_dumper_1877 = new("./chan_status1877.csv");
    fifo_monitor_1877 = new(fifo_csv_dumper_1877,fifo_intf_1877,cstatus_csv_dumper_1877);
    fifo_csv_dumper_1878 = new("./depth1878.csv");
    cstatus_csv_dumper_1878 = new("./chan_status1878.csv");
    fifo_monitor_1878 = new(fifo_csv_dumper_1878,fifo_intf_1878,cstatus_csv_dumper_1878);
    fifo_csv_dumper_1879 = new("./depth1879.csv");
    cstatus_csv_dumper_1879 = new("./chan_status1879.csv");
    fifo_monitor_1879 = new(fifo_csv_dumper_1879,fifo_intf_1879,cstatus_csv_dumper_1879);
    fifo_csv_dumper_1880 = new("./depth1880.csv");
    cstatus_csv_dumper_1880 = new("./chan_status1880.csv");
    fifo_monitor_1880 = new(fifo_csv_dumper_1880,fifo_intf_1880,cstatus_csv_dumper_1880);
    fifo_csv_dumper_1881 = new("./depth1881.csv");
    cstatus_csv_dumper_1881 = new("./chan_status1881.csv");
    fifo_monitor_1881 = new(fifo_csv_dumper_1881,fifo_intf_1881,cstatus_csv_dumper_1881);
    fifo_csv_dumper_1882 = new("./depth1882.csv");
    cstatus_csv_dumper_1882 = new("./chan_status1882.csv");
    fifo_monitor_1882 = new(fifo_csv_dumper_1882,fifo_intf_1882,cstatus_csv_dumper_1882);
    fifo_csv_dumper_1883 = new("./depth1883.csv");
    cstatus_csv_dumper_1883 = new("./chan_status1883.csv");
    fifo_monitor_1883 = new(fifo_csv_dumper_1883,fifo_intf_1883,cstatus_csv_dumper_1883);
    fifo_csv_dumper_1884 = new("./depth1884.csv");
    cstatus_csv_dumper_1884 = new("./chan_status1884.csv");
    fifo_monitor_1884 = new(fifo_csv_dumper_1884,fifo_intf_1884,cstatus_csv_dumper_1884);
    fifo_csv_dumper_1885 = new("./depth1885.csv");
    cstatus_csv_dumper_1885 = new("./chan_status1885.csv");
    fifo_monitor_1885 = new(fifo_csv_dumper_1885,fifo_intf_1885,cstatus_csv_dumper_1885);
    fifo_csv_dumper_1886 = new("./depth1886.csv");
    cstatus_csv_dumper_1886 = new("./chan_status1886.csv");
    fifo_monitor_1886 = new(fifo_csv_dumper_1886,fifo_intf_1886,cstatus_csv_dumper_1886);
    fifo_csv_dumper_1887 = new("./depth1887.csv");
    cstatus_csv_dumper_1887 = new("./chan_status1887.csv");
    fifo_monitor_1887 = new(fifo_csv_dumper_1887,fifo_intf_1887,cstatus_csv_dumper_1887);
    fifo_csv_dumper_1888 = new("./depth1888.csv");
    cstatus_csv_dumper_1888 = new("./chan_status1888.csv");
    fifo_monitor_1888 = new(fifo_csv_dumper_1888,fifo_intf_1888,cstatus_csv_dumper_1888);
    fifo_csv_dumper_1889 = new("./depth1889.csv");
    cstatus_csv_dumper_1889 = new("./chan_status1889.csv");
    fifo_monitor_1889 = new(fifo_csv_dumper_1889,fifo_intf_1889,cstatus_csv_dumper_1889);
    fifo_csv_dumper_1890 = new("./depth1890.csv");
    cstatus_csv_dumper_1890 = new("./chan_status1890.csv");
    fifo_monitor_1890 = new(fifo_csv_dumper_1890,fifo_intf_1890,cstatus_csv_dumper_1890);
    fifo_csv_dumper_1891 = new("./depth1891.csv");
    cstatus_csv_dumper_1891 = new("./chan_status1891.csv");
    fifo_monitor_1891 = new(fifo_csv_dumper_1891,fifo_intf_1891,cstatus_csv_dumper_1891);
    fifo_csv_dumper_1892 = new("./depth1892.csv");
    cstatus_csv_dumper_1892 = new("./chan_status1892.csv");
    fifo_monitor_1892 = new(fifo_csv_dumper_1892,fifo_intf_1892,cstatus_csv_dumper_1892);
    fifo_csv_dumper_1893 = new("./depth1893.csv");
    cstatus_csv_dumper_1893 = new("./chan_status1893.csv");
    fifo_monitor_1893 = new(fifo_csv_dumper_1893,fifo_intf_1893,cstatus_csv_dumper_1893);
    fifo_csv_dumper_1894 = new("./depth1894.csv");
    cstatus_csv_dumper_1894 = new("./chan_status1894.csv");
    fifo_monitor_1894 = new(fifo_csv_dumper_1894,fifo_intf_1894,cstatus_csv_dumper_1894);
    fifo_csv_dumper_1895 = new("./depth1895.csv");
    cstatus_csv_dumper_1895 = new("./chan_status1895.csv");
    fifo_monitor_1895 = new(fifo_csv_dumper_1895,fifo_intf_1895,cstatus_csv_dumper_1895);
    fifo_csv_dumper_1896 = new("./depth1896.csv");
    cstatus_csv_dumper_1896 = new("./chan_status1896.csv");
    fifo_monitor_1896 = new(fifo_csv_dumper_1896,fifo_intf_1896,cstatus_csv_dumper_1896);
    fifo_csv_dumper_1897 = new("./depth1897.csv");
    cstatus_csv_dumper_1897 = new("./chan_status1897.csv");
    fifo_monitor_1897 = new(fifo_csv_dumper_1897,fifo_intf_1897,cstatus_csv_dumper_1897);
    fifo_csv_dumper_1898 = new("./depth1898.csv");
    cstatus_csv_dumper_1898 = new("./chan_status1898.csv");
    fifo_monitor_1898 = new(fifo_csv_dumper_1898,fifo_intf_1898,cstatus_csv_dumper_1898);
    fifo_csv_dumper_1899 = new("./depth1899.csv");
    cstatus_csv_dumper_1899 = new("./chan_status1899.csv");
    fifo_monitor_1899 = new(fifo_csv_dumper_1899,fifo_intf_1899,cstatus_csv_dumper_1899);
    fifo_csv_dumper_1900 = new("./depth1900.csv");
    cstatus_csv_dumper_1900 = new("./chan_status1900.csv");
    fifo_monitor_1900 = new(fifo_csv_dumper_1900,fifo_intf_1900,cstatus_csv_dumper_1900);
    fifo_csv_dumper_1901 = new("./depth1901.csv");
    cstatus_csv_dumper_1901 = new("./chan_status1901.csv");
    fifo_monitor_1901 = new(fifo_csv_dumper_1901,fifo_intf_1901,cstatus_csv_dumper_1901);
    fifo_csv_dumper_1902 = new("./depth1902.csv");
    cstatus_csv_dumper_1902 = new("./chan_status1902.csv");
    fifo_monitor_1902 = new(fifo_csv_dumper_1902,fifo_intf_1902,cstatus_csv_dumper_1902);
    fifo_csv_dumper_1903 = new("./depth1903.csv");
    cstatus_csv_dumper_1903 = new("./chan_status1903.csv");
    fifo_monitor_1903 = new(fifo_csv_dumper_1903,fifo_intf_1903,cstatus_csv_dumper_1903);
    fifo_csv_dumper_1904 = new("./depth1904.csv");
    cstatus_csv_dumper_1904 = new("./chan_status1904.csv");
    fifo_monitor_1904 = new(fifo_csv_dumper_1904,fifo_intf_1904,cstatus_csv_dumper_1904);
    fifo_csv_dumper_1905 = new("./depth1905.csv");
    cstatus_csv_dumper_1905 = new("./chan_status1905.csv");
    fifo_monitor_1905 = new(fifo_csv_dumper_1905,fifo_intf_1905,cstatus_csv_dumper_1905);
    fifo_csv_dumper_1906 = new("./depth1906.csv");
    cstatus_csv_dumper_1906 = new("./chan_status1906.csv");
    fifo_monitor_1906 = new(fifo_csv_dumper_1906,fifo_intf_1906,cstatus_csv_dumper_1906);
    fifo_csv_dumper_1907 = new("./depth1907.csv");
    cstatus_csv_dumper_1907 = new("./chan_status1907.csv");
    fifo_monitor_1907 = new(fifo_csv_dumper_1907,fifo_intf_1907,cstatus_csv_dumper_1907);
    fifo_csv_dumper_1908 = new("./depth1908.csv");
    cstatus_csv_dumper_1908 = new("./chan_status1908.csv");
    fifo_monitor_1908 = new(fifo_csv_dumper_1908,fifo_intf_1908,cstatus_csv_dumper_1908);
    fifo_csv_dumper_1909 = new("./depth1909.csv");
    cstatus_csv_dumper_1909 = new("./chan_status1909.csv");
    fifo_monitor_1909 = new(fifo_csv_dumper_1909,fifo_intf_1909,cstatus_csv_dumper_1909);
    fifo_csv_dumper_1910 = new("./depth1910.csv");
    cstatus_csv_dumper_1910 = new("./chan_status1910.csv");
    fifo_monitor_1910 = new(fifo_csv_dumper_1910,fifo_intf_1910,cstatus_csv_dumper_1910);
    fifo_csv_dumper_1911 = new("./depth1911.csv");
    cstatus_csv_dumper_1911 = new("./chan_status1911.csv");
    fifo_monitor_1911 = new(fifo_csv_dumper_1911,fifo_intf_1911,cstatus_csv_dumper_1911);
    fifo_csv_dumper_1912 = new("./depth1912.csv");
    cstatus_csv_dumper_1912 = new("./chan_status1912.csv");
    fifo_monitor_1912 = new(fifo_csv_dumper_1912,fifo_intf_1912,cstatus_csv_dumper_1912);
    fifo_csv_dumper_1913 = new("./depth1913.csv");
    cstatus_csv_dumper_1913 = new("./chan_status1913.csv");
    fifo_monitor_1913 = new(fifo_csv_dumper_1913,fifo_intf_1913,cstatus_csv_dumper_1913);
    fifo_csv_dumper_1914 = new("./depth1914.csv");
    cstatus_csv_dumper_1914 = new("./chan_status1914.csv");
    fifo_monitor_1914 = new(fifo_csv_dumper_1914,fifo_intf_1914,cstatus_csv_dumper_1914);
    fifo_csv_dumper_1915 = new("./depth1915.csv");
    cstatus_csv_dumper_1915 = new("./chan_status1915.csv");
    fifo_monitor_1915 = new(fifo_csv_dumper_1915,fifo_intf_1915,cstatus_csv_dumper_1915);
    fifo_csv_dumper_1916 = new("./depth1916.csv");
    cstatus_csv_dumper_1916 = new("./chan_status1916.csv");
    fifo_monitor_1916 = new(fifo_csv_dumper_1916,fifo_intf_1916,cstatus_csv_dumper_1916);
    fifo_csv_dumper_1917 = new("./depth1917.csv");
    cstatus_csv_dumper_1917 = new("./chan_status1917.csv");
    fifo_monitor_1917 = new(fifo_csv_dumper_1917,fifo_intf_1917,cstatus_csv_dumper_1917);
    fifo_csv_dumper_1918 = new("./depth1918.csv");
    cstatus_csv_dumper_1918 = new("./chan_status1918.csv");
    fifo_monitor_1918 = new(fifo_csv_dumper_1918,fifo_intf_1918,cstatus_csv_dumper_1918);
    fifo_csv_dumper_1919 = new("./depth1919.csv");
    cstatus_csv_dumper_1919 = new("./chan_status1919.csv");
    fifo_monitor_1919 = new(fifo_csv_dumper_1919,fifo_intf_1919,cstatus_csv_dumper_1919);
    fifo_csv_dumper_1920 = new("./depth1920.csv");
    cstatus_csv_dumper_1920 = new("./chan_status1920.csv");
    fifo_monitor_1920 = new(fifo_csv_dumper_1920,fifo_intf_1920,cstatus_csv_dumper_1920);
    fifo_csv_dumper_1921 = new("./depth1921.csv");
    cstatus_csv_dumper_1921 = new("./chan_status1921.csv");
    fifo_monitor_1921 = new(fifo_csv_dumper_1921,fifo_intf_1921,cstatus_csv_dumper_1921);
    fifo_csv_dumper_1922 = new("./depth1922.csv");
    cstatus_csv_dumper_1922 = new("./chan_status1922.csv");
    fifo_monitor_1922 = new(fifo_csv_dumper_1922,fifo_intf_1922,cstatus_csv_dumper_1922);
    fifo_csv_dumper_1923 = new("./depth1923.csv");
    cstatus_csv_dumper_1923 = new("./chan_status1923.csv");
    fifo_monitor_1923 = new(fifo_csv_dumper_1923,fifo_intf_1923,cstatus_csv_dumper_1923);
    fifo_csv_dumper_1924 = new("./depth1924.csv");
    cstatus_csv_dumper_1924 = new("./chan_status1924.csv");
    fifo_monitor_1924 = new(fifo_csv_dumper_1924,fifo_intf_1924,cstatus_csv_dumper_1924);
    fifo_csv_dumper_1925 = new("./depth1925.csv");
    cstatus_csv_dumper_1925 = new("./chan_status1925.csv");
    fifo_monitor_1925 = new(fifo_csv_dumper_1925,fifo_intf_1925,cstatus_csv_dumper_1925);
    fifo_csv_dumper_1926 = new("./depth1926.csv");
    cstatus_csv_dumper_1926 = new("./chan_status1926.csv");
    fifo_monitor_1926 = new(fifo_csv_dumper_1926,fifo_intf_1926,cstatus_csv_dumper_1926);
    fifo_csv_dumper_1927 = new("./depth1927.csv");
    cstatus_csv_dumper_1927 = new("./chan_status1927.csv");
    fifo_monitor_1927 = new(fifo_csv_dumper_1927,fifo_intf_1927,cstatus_csv_dumper_1927);
    fifo_csv_dumper_1928 = new("./depth1928.csv");
    cstatus_csv_dumper_1928 = new("./chan_status1928.csv");
    fifo_monitor_1928 = new(fifo_csv_dumper_1928,fifo_intf_1928,cstatus_csv_dumper_1928);
    fifo_csv_dumper_1929 = new("./depth1929.csv");
    cstatus_csv_dumper_1929 = new("./chan_status1929.csv");
    fifo_monitor_1929 = new(fifo_csv_dumper_1929,fifo_intf_1929,cstatus_csv_dumper_1929);
    fifo_csv_dumper_1930 = new("./depth1930.csv");
    cstatus_csv_dumper_1930 = new("./chan_status1930.csv");
    fifo_monitor_1930 = new(fifo_csv_dumper_1930,fifo_intf_1930,cstatus_csv_dumper_1930);
    fifo_csv_dumper_1931 = new("./depth1931.csv");
    cstatus_csv_dumper_1931 = new("./chan_status1931.csv");
    fifo_monitor_1931 = new(fifo_csv_dumper_1931,fifo_intf_1931,cstatus_csv_dumper_1931);
    fifo_csv_dumper_1932 = new("./depth1932.csv");
    cstatus_csv_dumper_1932 = new("./chan_status1932.csv");
    fifo_monitor_1932 = new(fifo_csv_dumper_1932,fifo_intf_1932,cstatus_csv_dumper_1932);
    fifo_csv_dumper_1933 = new("./depth1933.csv");
    cstatus_csv_dumper_1933 = new("./chan_status1933.csv");
    fifo_monitor_1933 = new(fifo_csv_dumper_1933,fifo_intf_1933,cstatus_csv_dumper_1933);
    fifo_csv_dumper_1934 = new("./depth1934.csv");
    cstatus_csv_dumper_1934 = new("./chan_status1934.csv");
    fifo_monitor_1934 = new(fifo_csv_dumper_1934,fifo_intf_1934,cstatus_csv_dumper_1934);
    fifo_csv_dumper_1935 = new("./depth1935.csv");
    cstatus_csv_dumper_1935 = new("./chan_status1935.csv");
    fifo_monitor_1935 = new(fifo_csv_dumper_1935,fifo_intf_1935,cstatus_csv_dumper_1935);
    fifo_csv_dumper_1936 = new("./depth1936.csv");
    cstatus_csv_dumper_1936 = new("./chan_status1936.csv");
    fifo_monitor_1936 = new(fifo_csv_dumper_1936,fifo_intf_1936,cstatus_csv_dumper_1936);
    fifo_csv_dumper_1937 = new("./depth1937.csv");
    cstatus_csv_dumper_1937 = new("./chan_status1937.csv");
    fifo_monitor_1937 = new(fifo_csv_dumper_1937,fifo_intf_1937,cstatus_csv_dumper_1937);
    fifo_csv_dumper_1938 = new("./depth1938.csv");
    cstatus_csv_dumper_1938 = new("./chan_status1938.csv");
    fifo_monitor_1938 = new(fifo_csv_dumper_1938,fifo_intf_1938,cstatus_csv_dumper_1938);
    fifo_csv_dumper_1939 = new("./depth1939.csv");
    cstatus_csv_dumper_1939 = new("./chan_status1939.csv");
    fifo_monitor_1939 = new(fifo_csv_dumper_1939,fifo_intf_1939,cstatus_csv_dumper_1939);
    fifo_csv_dumper_1940 = new("./depth1940.csv");
    cstatus_csv_dumper_1940 = new("./chan_status1940.csv");
    fifo_monitor_1940 = new(fifo_csv_dumper_1940,fifo_intf_1940,cstatus_csv_dumper_1940);
    fifo_csv_dumper_1941 = new("./depth1941.csv");
    cstatus_csv_dumper_1941 = new("./chan_status1941.csv");
    fifo_monitor_1941 = new(fifo_csv_dumper_1941,fifo_intf_1941,cstatus_csv_dumper_1941);
    fifo_csv_dumper_1942 = new("./depth1942.csv");
    cstatus_csv_dumper_1942 = new("./chan_status1942.csv");
    fifo_monitor_1942 = new(fifo_csv_dumper_1942,fifo_intf_1942,cstatus_csv_dumper_1942);
    fifo_csv_dumper_1943 = new("./depth1943.csv");
    cstatus_csv_dumper_1943 = new("./chan_status1943.csv");
    fifo_monitor_1943 = new(fifo_csv_dumper_1943,fifo_intf_1943,cstatus_csv_dumper_1943);
    fifo_csv_dumper_1944 = new("./depth1944.csv");
    cstatus_csv_dumper_1944 = new("./chan_status1944.csv");
    fifo_monitor_1944 = new(fifo_csv_dumper_1944,fifo_intf_1944,cstatus_csv_dumper_1944);
    fifo_csv_dumper_1945 = new("./depth1945.csv");
    cstatus_csv_dumper_1945 = new("./chan_status1945.csv");
    fifo_monitor_1945 = new(fifo_csv_dumper_1945,fifo_intf_1945,cstatus_csv_dumper_1945);
    fifo_csv_dumper_1946 = new("./depth1946.csv");
    cstatus_csv_dumper_1946 = new("./chan_status1946.csv");
    fifo_monitor_1946 = new(fifo_csv_dumper_1946,fifo_intf_1946,cstatus_csv_dumper_1946);
    fifo_csv_dumper_1947 = new("./depth1947.csv");
    cstatus_csv_dumper_1947 = new("./chan_status1947.csv");
    fifo_monitor_1947 = new(fifo_csv_dumper_1947,fifo_intf_1947,cstatus_csv_dumper_1947);
    fifo_csv_dumper_1948 = new("./depth1948.csv");
    cstatus_csv_dumper_1948 = new("./chan_status1948.csv");
    fifo_monitor_1948 = new(fifo_csv_dumper_1948,fifo_intf_1948,cstatus_csv_dumper_1948);
    fifo_csv_dumper_1949 = new("./depth1949.csv");
    cstatus_csv_dumper_1949 = new("./chan_status1949.csv");
    fifo_monitor_1949 = new(fifo_csv_dumper_1949,fifo_intf_1949,cstatus_csv_dumper_1949);
    fifo_csv_dumper_1950 = new("./depth1950.csv");
    cstatus_csv_dumper_1950 = new("./chan_status1950.csv");
    fifo_monitor_1950 = new(fifo_csv_dumper_1950,fifo_intf_1950,cstatus_csv_dumper_1950);
    fifo_csv_dumper_1951 = new("./depth1951.csv");
    cstatus_csv_dumper_1951 = new("./chan_status1951.csv");
    fifo_monitor_1951 = new(fifo_csv_dumper_1951,fifo_intf_1951,cstatus_csv_dumper_1951);
    fifo_csv_dumper_1952 = new("./depth1952.csv");
    cstatus_csv_dumper_1952 = new("./chan_status1952.csv");
    fifo_monitor_1952 = new(fifo_csv_dumper_1952,fifo_intf_1952,cstatus_csv_dumper_1952);
    fifo_csv_dumper_1953 = new("./depth1953.csv");
    cstatus_csv_dumper_1953 = new("./chan_status1953.csv");
    fifo_monitor_1953 = new(fifo_csv_dumper_1953,fifo_intf_1953,cstatus_csv_dumper_1953);
    fifo_csv_dumper_1954 = new("./depth1954.csv");
    cstatus_csv_dumper_1954 = new("./chan_status1954.csv");
    fifo_monitor_1954 = new(fifo_csv_dumper_1954,fifo_intf_1954,cstatus_csv_dumper_1954);
    fifo_csv_dumper_1955 = new("./depth1955.csv");
    cstatus_csv_dumper_1955 = new("./chan_status1955.csv");
    fifo_monitor_1955 = new(fifo_csv_dumper_1955,fifo_intf_1955,cstatus_csv_dumper_1955);
    fifo_csv_dumper_1956 = new("./depth1956.csv");
    cstatus_csv_dumper_1956 = new("./chan_status1956.csv");
    fifo_monitor_1956 = new(fifo_csv_dumper_1956,fifo_intf_1956,cstatus_csv_dumper_1956);
    fifo_csv_dumper_1957 = new("./depth1957.csv");
    cstatus_csv_dumper_1957 = new("./chan_status1957.csv");
    fifo_monitor_1957 = new(fifo_csv_dumper_1957,fifo_intf_1957,cstatus_csv_dumper_1957);
    fifo_csv_dumper_1958 = new("./depth1958.csv");
    cstatus_csv_dumper_1958 = new("./chan_status1958.csv");
    fifo_monitor_1958 = new(fifo_csv_dumper_1958,fifo_intf_1958,cstatus_csv_dumper_1958);
    fifo_csv_dumper_1959 = new("./depth1959.csv");
    cstatus_csv_dumper_1959 = new("./chan_status1959.csv");
    fifo_monitor_1959 = new(fifo_csv_dumper_1959,fifo_intf_1959,cstatus_csv_dumper_1959);
    fifo_csv_dumper_1960 = new("./depth1960.csv");
    cstatus_csv_dumper_1960 = new("./chan_status1960.csv");
    fifo_monitor_1960 = new(fifo_csv_dumper_1960,fifo_intf_1960,cstatus_csv_dumper_1960);
    fifo_csv_dumper_1961 = new("./depth1961.csv");
    cstatus_csv_dumper_1961 = new("./chan_status1961.csv");
    fifo_monitor_1961 = new(fifo_csv_dumper_1961,fifo_intf_1961,cstatus_csv_dumper_1961);
    fifo_csv_dumper_1962 = new("./depth1962.csv");
    cstatus_csv_dumper_1962 = new("./chan_status1962.csv");
    fifo_monitor_1962 = new(fifo_csv_dumper_1962,fifo_intf_1962,cstatus_csv_dumper_1962);
    fifo_csv_dumper_1963 = new("./depth1963.csv");
    cstatus_csv_dumper_1963 = new("./chan_status1963.csv");
    fifo_monitor_1963 = new(fifo_csv_dumper_1963,fifo_intf_1963,cstatus_csv_dumper_1963);
    fifo_csv_dumper_1964 = new("./depth1964.csv");
    cstatus_csv_dumper_1964 = new("./chan_status1964.csv");
    fifo_monitor_1964 = new(fifo_csv_dumper_1964,fifo_intf_1964,cstatus_csv_dumper_1964);
    fifo_csv_dumper_1965 = new("./depth1965.csv");
    cstatus_csv_dumper_1965 = new("./chan_status1965.csv");
    fifo_monitor_1965 = new(fifo_csv_dumper_1965,fifo_intf_1965,cstatus_csv_dumper_1965);
    fifo_csv_dumper_1966 = new("./depth1966.csv");
    cstatus_csv_dumper_1966 = new("./chan_status1966.csv");
    fifo_monitor_1966 = new(fifo_csv_dumper_1966,fifo_intf_1966,cstatus_csv_dumper_1966);
    fifo_csv_dumper_1967 = new("./depth1967.csv");
    cstatus_csv_dumper_1967 = new("./chan_status1967.csv");
    fifo_monitor_1967 = new(fifo_csv_dumper_1967,fifo_intf_1967,cstatus_csv_dumper_1967);
    fifo_csv_dumper_1968 = new("./depth1968.csv");
    cstatus_csv_dumper_1968 = new("./chan_status1968.csv");
    fifo_monitor_1968 = new(fifo_csv_dumper_1968,fifo_intf_1968,cstatus_csv_dumper_1968);
    fifo_csv_dumper_1969 = new("./depth1969.csv");
    cstatus_csv_dumper_1969 = new("./chan_status1969.csv");
    fifo_monitor_1969 = new(fifo_csv_dumper_1969,fifo_intf_1969,cstatus_csv_dumper_1969);
    fifo_csv_dumper_1970 = new("./depth1970.csv");
    cstatus_csv_dumper_1970 = new("./chan_status1970.csv");
    fifo_monitor_1970 = new(fifo_csv_dumper_1970,fifo_intf_1970,cstatus_csv_dumper_1970);
    fifo_csv_dumper_1971 = new("./depth1971.csv");
    cstatus_csv_dumper_1971 = new("./chan_status1971.csv");
    fifo_monitor_1971 = new(fifo_csv_dumper_1971,fifo_intf_1971,cstatus_csv_dumper_1971);
    fifo_csv_dumper_1972 = new("./depth1972.csv");
    cstatus_csv_dumper_1972 = new("./chan_status1972.csv");
    fifo_monitor_1972 = new(fifo_csv_dumper_1972,fifo_intf_1972,cstatus_csv_dumper_1972);
    fifo_csv_dumper_1973 = new("./depth1973.csv");
    cstatus_csv_dumper_1973 = new("./chan_status1973.csv");
    fifo_monitor_1973 = new(fifo_csv_dumper_1973,fifo_intf_1973,cstatus_csv_dumper_1973);
    fifo_csv_dumper_1974 = new("./depth1974.csv");
    cstatus_csv_dumper_1974 = new("./chan_status1974.csv");
    fifo_monitor_1974 = new(fifo_csv_dumper_1974,fifo_intf_1974,cstatus_csv_dumper_1974);
    fifo_csv_dumper_1975 = new("./depth1975.csv");
    cstatus_csv_dumper_1975 = new("./chan_status1975.csv");
    fifo_monitor_1975 = new(fifo_csv_dumper_1975,fifo_intf_1975,cstatus_csv_dumper_1975);
    fifo_csv_dumper_1976 = new("./depth1976.csv");
    cstatus_csv_dumper_1976 = new("./chan_status1976.csv");
    fifo_monitor_1976 = new(fifo_csv_dumper_1976,fifo_intf_1976,cstatus_csv_dumper_1976);
    fifo_csv_dumper_1977 = new("./depth1977.csv");
    cstatus_csv_dumper_1977 = new("./chan_status1977.csv");
    fifo_monitor_1977 = new(fifo_csv_dumper_1977,fifo_intf_1977,cstatus_csv_dumper_1977);
    fifo_csv_dumper_1978 = new("./depth1978.csv");
    cstatus_csv_dumper_1978 = new("./chan_status1978.csv");
    fifo_monitor_1978 = new(fifo_csv_dumper_1978,fifo_intf_1978,cstatus_csv_dumper_1978);
    fifo_csv_dumper_1979 = new("./depth1979.csv");
    cstatus_csv_dumper_1979 = new("./chan_status1979.csv");
    fifo_monitor_1979 = new(fifo_csv_dumper_1979,fifo_intf_1979,cstatus_csv_dumper_1979);
    fifo_csv_dumper_1980 = new("./depth1980.csv");
    cstatus_csv_dumper_1980 = new("./chan_status1980.csv");
    fifo_monitor_1980 = new(fifo_csv_dumper_1980,fifo_intf_1980,cstatus_csv_dumper_1980);
    fifo_csv_dumper_1981 = new("./depth1981.csv");
    cstatus_csv_dumper_1981 = new("./chan_status1981.csv");
    fifo_monitor_1981 = new(fifo_csv_dumper_1981,fifo_intf_1981,cstatus_csv_dumper_1981);
    fifo_csv_dumper_1982 = new("./depth1982.csv");
    cstatus_csv_dumper_1982 = new("./chan_status1982.csv");
    fifo_monitor_1982 = new(fifo_csv_dumper_1982,fifo_intf_1982,cstatus_csv_dumper_1982);
    fifo_csv_dumper_1983 = new("./depth1983.csv");
    cstatus_csv_dumper_1983 = new("./chan_status1983.csv");
    fifo_monitor_1983 = new(fifo_csv_dumper_1983,fifo_intf_1983,cstatus_csv_dumper_1983);
    fifo_csv_dumper_1984 = new("./depth1984.csv");
    cstatus_csv_dumper_1984 = new("./chan_status1984.csv");
    fifo_monitor_1984 = new(fifo_csv_dumper_1984,fifo_intf_1984,cstatus_csv_dumper_1984);
    fifo_csv_dumper_1985 = new("./depth1985.csv");
    cstatus_csv_dumper_1985 = new("./chan_status1985.csv");
    fifo_monitor_1985 = new(fifo_csv_dumper_1985,fifo_intf_1985,cstatus_csv_dumper_1985);
    fifo_csv_dumper_1986 = new("./depth1986.csv");
    cstatus_csv_dumper_1986 = new("./chan_status1986.csv");
    fifo_monitor_1986 = new(fifo_csv_dumper_1986,fifo_intf_1986,cstatus_csv_dumper_1986);
    fifo_csv_dumper_1987 = new("./depth1987.csv");
    cstatus_csv_dumper_1987 = new("./chan_status1987.csv");
    fifo_monitor_1987 = new(fifo_csv_dumper_1987,fifo_intf_1987,cstatus_csv_dumper_1987);
    fifo_csv_dumper_1988 = new("./depth1988.csv");
    cstatus_csv_dumper_1988 = new("./chan_status1988.csv");
    fifo_monitor_1988 = new(fifo_csv_dumper_1988,fifo_intf_1988,cstatus_csv_dumper_1988);
    fifo_csv_dumper_1989 = new("./depth1989.csv");
    cstatus_csv_dumper_1989 = new("./chan_status1989.csv");
    fifo_monitor_1989 = new(fifo_csv_dumper_1989,fifo_intf_1989,cstatus_csv_dumper_1989);
    fifo_csv_dumper_1990 = new("./depth1990.csv");
    cstatus_csv_dumper_1990 = new("./chan_status1990.csv");
    fifo_monitor_1990 = new(fifo_csv_dumper_1990,fifo_intf_1990,cstatus_csv_dumper_1990);
    fifo_csv_dumper_1991 = new("./depth1991.csv");
    cstatus_csv_dumper_1991 = new("./chan_status1991.csv");
    fifo_monitor_1991 = new(fifo_csv_dumper_1991,fifo_intf_1991,cstatus_csv_dumper_1991);
    fifo_csv_dumper_1992 = new("./depth1992.csv");
    cstatus_csv_dumper_1992 = new("./chan_status1992.csv");
    fifo_monitor_1992 = new(fifo_csv_dumper_1992,fifo_intf_1992,cstatus_csv_dumper_1992);
    fifo_csv_dumper_1993 = new("./depth1993.csv");
    cstatus_csv_dumper_1993 = new("./chan_status1993.csv");
    fifo_monitor_1993 = new(fifo_csv_dumper_1993,fifo_intf_1993,cstatus_csv_dumper_1993);
    fifo_csv_dumper_1994 = new("./depth1994.csv");
    cstatus_csv_dumper_1994 = new("./chan_status1994.csv");
    fifo_monitor_1994 = new(fifo_csv_dumper_1994,fifo_intf_1994,cstatus_csv_dumper_1994);
    fifo_csv_dumper_1995 = new("./depth1995.csv");
    cstatus_csv_dumper_1995 = new("./chan_status1995.csv");
    fifo_monitor_1995 = new(fifo_csv_dumper_1995,fifo_intf_1995,cstatus_csv_dumper_1995);
    fifo_csv_dumper_1996 = new("./depth1996.csv");
    cstatus_csv_dumper_1996 = new("./chan_status1996.csv");
    fifo_monitor_1996 = new(fifo_csv_dumper_1996,fifo_intf_1996,cstatus_csv_dumper_1996);
    fifo_csv_dumper_1997 = new("./depth1997.csv");
    cstatus_csv_dumper_1997 = new("./chan_status1997.csv");
    fifo_monitor_1997 = new(fifo_csv_dumper_1997,fifo_intf_1997,cstatus_csv_dumper_1997);
    fifo_csv_dumper_1998 = new("./depth1998.csv");
    cstatus_csv_dumper_1998 = new("./chan_status1998.csv");
    fifo_monitor_1998 = new(fifo_csv_dumper_1998,fifo_intf_1998,cstatus_csv_dumper_1998);
    fifo_csv_dumper_1999 = new("./depth1999.csv");
    cstatus_csv_dumper_1999 = new("./chan_status1999.csv");
    fifo_monitor_1999 = new(fifo_csv_dumper_1999,fifo_intf_1999,cstatus_csv_dumper_1999);
    fifo_csv_dumper_2000 = new("./depth2000.csv");
    cstatus_csv_dumper_2000 = new("./chan_status2000.csv");
    fifo_monitor_2000 = new(fifo_csv_dumper_2000,fifo_intf_2000,cstatus_csv_dumper_2000);
    fifo_csv_dumper_2001 = new("./depth2001.csv");
    cstatus_csv_dumper_2001 = new("./chan_status2001.csv");
    fifo_monitor_2001 = new(fifo_csv_dumper_2001,fifo_intf_2001,cstatus_csv_dumper_2001);
    fifo_csv_dumper_2002 = new("./depth2002.csv");
    cstatus_csv_dumper_2002 = new("./chan_status2002.csv");
    fifo_monitor_2002 = new(fifo_csv_dumper_2002,fifo_intf_2002,cstatus_csv_dumper_2002);
    fifo_csv_dumper_2003 = new("./depth2003.csv");
    cstatus_csv_dumper_2003 = new("./chan_status2003.csv");
    fifo_monitor_2003 = new(fifo_csv_dumper_2003,fifo_intf_2003,cstatus_csv_dumper_2003);
    fifo_csv_dumper_2004 = new("./depth2004.csv");
    cstatus_csv_dumper_2004 = new("./chan_status2004.csv");
    fifo_monitor_2004 = new(fifo_csv_dumper_2004,fifo_intf_2004,cstatus_csv_dumper_2004);
    fifo_csv_dumper_2005 = new("./depth2005.csv");
    cstatus_csv_dumper_2005 = new("./chan_status2005.csv");
    fifo_monitor_2005 = new(fifo_csv_dumper_2005,fifo_intf_2005,cstatus_csv_dumper_2005);
    fifo_csv_dumper_2006 = new("./depth2006.csv");
    cstatus_csv_dumper_2006 = new("./chan_status2006.csv");
    fifo_monitor_2006 = new(fifo_csv_dumper_2006,fifo_intf_2006,cstatus_csv_dumper_2006);
    fifo_csv_dumper_2007 = new("./depth2007.csv");
    cstatus_csv_dumper_2007 = new("./chan_status2007.csv");
    fifo_monitor_2007 = new(fifo_csv_dumper_2007,fifo_intf_2007,cstatus_csv_dumper_2007);
    fifo_csv_dumper_2008 = new("./depth2008.csv");
    cstatus_csv_dumper_2008 = new("./chan_status2008.csv");
    fifo_monitor_2008 = new(fifo_csv_dumper_2008,fifo_intf_2008,cstatus_csv_dumper_2008);
    fifo_csv_dumper_2009 = new("./depth2009.csv");
    cstatus_csv_dumper_2009 = new("./chan_status2009.csv");
    fifo_monitor_2009 = new(fifo_csv_dumper_2009,fifo_intf_2009,cstatus_csv_dumper_2009);
    fifo_csv_dumper_2010 = new("./depth2010.csv");
    cstatus_csv_dumper_2010 = new("./chan_status2010.csv");
    fifo_monitor_2010 = new(fifo_csv_dumper_2010,fifo_intf_2010,cstatus_csv_dumper_2010);
    fifo_csv_dumper_2011 = new("./depth2011.csv");
    cstatus_csv_dumper_2011 = new("./chan_status2011.csv");
    fifo_monitor_2011 = new(fifo_csv_dumper_2011,fifo_intf_2011,cstatus_csv_dumper_2011);
    fifo_csv_dumper_2012 = new("./depth2012.csv");
    cstatus_csv_dumper_2012 = new("./chan_status2012.csv");
    fifo_monitor_2012 = new(fifo_csv_dumper_2012,fifo_intf_2012,cstatus_csv_dumper_2012);
    fifo_csv_dumper_2013 = new("./depth2013.csv");
    cstatus_csv_dumper_2013 = new("./chan_status2013.csv");
    fifo_monitor_2013 = new(fifo_csv_dumper_2013,fifo_intf_2013,cstatus_csv_dumper_2013);
    fifo_csv_dumper_2014 = new("./depth2014.csv");
    cstatus_csv_dumper_2014 = new("./chan_status2014.csv");
    fifo_monitor_2014 = new(fifo_csv_dumper_2014,fifo_intf_2014,cstatus_csv_dumper_2014);
    fifo_csv_dumper_2015 = new("./depth2015.csv");
    cstatus_csv_dumper_2015 = new("./chan_status2015.csv");
    fifo_monitor_2015 = new(fifo_csv_dumper_2015,fifo_intf_2015,cstatus_csv_dumper_2015);
    fifo_csv_dumper_2016 = new("./depth2016.csv");
    cstatus_csv_dumper_2016 = new("./chan_status2016.csv");
    fifo_monitor_2016 = new(fifo_csv_dumper_2016,fifo_intf_2016,cstatus_csv_dumper_2016);
    fifo_csv_dumper_2017 = new("./depth2017.csv");
    cstatus_csv_dumper_2017 = new("./chan_status2017.csv");
    fifo_monitor_2017 = new(fifo_csv_dumper_2017,fifo_intf_2017,cstatus_csv_dumper_2017);
    fifo_csv_dumper_2018 = new("./depth2018.csv");
    cstatus_csv_dumper_2018 = new("./chan_status2018.csv");
    fifo_monitor_2018 = new(fifo_csv_dumper_2018,fifo_intf_2018,cstatus_csv_dumper_2018);
    fifo_csv_dumper_2019 = new("./depth2019.csv");
    cstatus_csv_dumper_2019 = new("./chan_status2019.csv");
    fifo_monitor_2019 = new(fifo_csv_dumper_2019,fifo_intf_2019,cstatus_csv_dumper_2019);
    fifo_csv_dumper_2020 = new("./depth2020.csv");
    cstatus_csv_dumper_2020 = new("./chan_status2020.csv");
    fifo_monitor_2020 = new(fifo_csv_dumper_2020,fifo_intf_2020,cstatus_csv_dumper_2020);
    fifo_csv_dumper_2021 = new("./depth2021.csv");
    cstatus_csv_dumper_2021 = new("./chan_status2021.csv");
    fifo_monitor_2021 = new(fifo_csv_dumper_2021,fifo_intf_2021,cstatus_csv_dumper_2021);
    fifo_csv_dumper_2022 = new("./depth2022.csv");
    cstatus_csv_dumper_2022 = new("./chan_status2022.csv");
    fifo_monitor_2022 = new(fifo_csv_dumper_2022,fifo_intf_2022,cstatus_csv_dumper_2022);
    fifo_csv_dumper_2023 = new("./depth2023.csv");
    cstatus_csv_dumper_2023 = new("./chan_status2023.csv");
    fifo_monitor_2023 = new(fifo_csv_dumper_2023,fifo_intf_2023,cstatus_csv_dumper_2023);
    fifo_csv_dumper_2024 = new("./depth2024.csv");
    cstatus_csv_dumper_2024 = new("./chan_status2024.csv");
    fifo_monitor_2024 = new(fifo_csv_dumper_2024,fifo_intf_2024,cstatus_csv_dumper_2024);
    fifo_csv_dumper_2025 = new("./depth2025.csv");
    cstatus_csv_dumper_2025 = new("./chan_status2025.csv");
    fifo_monitor_2025 = new(fifo_csv_dumper_2025,fifo_intf_2025,cstatus_csv_dumper_2025);
    fifo_csv_dumper_2026 = new("./depth2026.csv");
    cstatus_csv_dumper_2026 = new("./chan_status2026.csv");
    fifo_monitor_2026 = new(fifo_csv_dumper_2026,fifo_intf_2026,cstatus_csv_dumper_2026);
    fifo_csv_dumper_2027 = new("./depth2027.csv");
    cstatus_csv_dumper_2027 = new("./chan_status2027.csv");
    fifo_monitor_2027 = new(fifo_csv_dumper_2027,fifo_intf_2027,cstatus_csv_dumper_2027);
    fifo_csv_dumper_2028 = new("./depth2028.csv");
    cstatus_csv_dumper_2028 = new("./chan_status2028.csv");
    fifo_monitor_2028 = new(fifo_csv_dumper_2028,fifo_intf_2028,cstatus_csv_dumper_2028);
    fifo_csv_dumper_2029 = new("./depth2029.csv");
    cstatus_csv_dumper_2029 = new("./chan_status2029.csv");
    fifo_monitor_2029 = new(fifo_csv_dumper_2029,fifo_intf_2029,cstatus_csv_dumper_2029);
    fifo_csv_dumper_2030 = new("./depth2030.csv");
    cstatus_csv_dumper_2030 = new("./chan_status2030.csv");
    fifo_monitor_2030 = new(fifo_csv_dumper_2030,fifo_intf_2030,cstatus_csv_dumper_2030);
    fifo_csv_dumper_2031 = new("./depth2031.csv");
    cstatus_csv_dumper_2031 = new("./chan_status2031.csv");
    fifo_monitor_2031 = new(fifo_csv_dumper_2031,fifo_intf_2031,cstatus_csv_dumper_2031);
    fifo_csv_dumper_2032 = new("./depth2032.csv");
    cstatus_csv_dumper_2032 = new("./chan_status2032.csv");
    fifo_monitor_2032 = new(fifo_csv_dumper_2032,fifo_intf_2032,cstatus_csv_dumper_2032);
    fifo_csv_dumper_2033 = new("./depth2033.csv");
    cstatus_csv_dumper_2033 = new("./chan_status2033.csv");
    fifo_monitor_2033 = new(fifo_csv_dumper_2033,fifo_intf_2033,cstatus_csv_dumper_2033);
    fifo_csv_dumper_2034 = new("./depth2034.csv");
    cstatus_csv_dumper_2034 = new("./chan_status2034.csv");
    fifo_monitor_2034 = new(fifo_csv_dumper_2034,fifo_intf_2034,cstatus_csv_dumper_2034);
    fifo_csv_dumper_2035 = new("./depth2035.csv");
    cstatus_csv_dumper_2035 = new("./chan_status2035.csv");
    fifo_monitor_2035 = new(fifo_csv_dumper_2035,fifo_intf_2035,cstatus_csv_dumper_2035);
    fifo_csv_dumper_2036 = new("./depth2036.csv");
    cstatus_csv_dumper_2036 = new("./chan_status2036.csv");
    fifo_monitor_2036 = new(fifo_csv_dumper_2036,fifo_intf_2036,cstatus_csv_dumper_2036);
    fifo_csv_dumper_2037 = new("./depth2037.csv");
    cstatus_csv_dumper_2037 = new("./chan_status2037.csv");
    fifo_monitor_2037 = new(fifo_csv_dumper_2037,fifo_intf_2037,cstatus_csv_dumper_2037);
    fifo_csv_dumper_2038 = new("./depth2038.csv");
    cstatus_csv_dumper_2038 = new("./chan_status2038.csv");
    fifo_monitor_2038 = new(fifo_csv_dumper_2038,fifo_intf_2038,cstatus_csv_dumper_2038);
    fifo_csv_dumper_2039 = new("./depth2039.csv");
    cstatus_csv_dumper_2039 = new("./chan_status2039.csv");
    fifo_monitor_2039 = new(fifo_csv_dumper_2039,fifo_intf_2039,cstatus_csv_dumper_2039);
    fifo_csv_dumper_2040 = new("./depth2040.csv");
    cstatus_csv_dumper_2040 = new("./chan_status2040.csv");
    fifo_monitor_2040 = new(fifo_csv_dumper_2040,fifo_intf_2040,cstatus_csv_dumper_2040);
    fifo_csv_dumper_2041 = new("./depth2041.csv");
    cstatus_csv_dumper_2041 = new("./chan_status2041.csv");
    fifo_monitor_2041 = new(fifo_csv_dumper_2041,fifo_intf_2041,cstatus_csv_dumper_2041);
    fifo_csv_dumper_2042 = new("./depth2042.csv");
    cstatus_csv_dumper_2042 = new("./chan_status2042.csv");
    fifo_monitor_2042 = new(fifo_csv_dumper_2042,fifo_intf_2042,cstatus_csv_dumper_2042);
    fifo_csv_dumper_2043 = new("./depth2043.csv");
    cstatus_csv_dumper_2043 = new("./chan_status2043.csv");
    fifo_monitor_2043 = new(fifo_csv_dumper_2043,fifo_intf_2043,cstatus_csv_dumper_2043);
    fifo_csv_dumper_2044 = new("./depth2044.csv");
    cstatus_csv_dumper_2044 = new("./chan_status2044.csv");
    fifo_monitor_2044 = new(fifo_csv_dumper_2044,fifo_intf_2044,cstatus_csv_dumper_2044);
    fifo_csv_dumper_2045 = new("./depth2045.csv");
    cstatus_csv_dumper_2045 = new("./chan_status2045.csv");
    fifo_monitor_2045 = new(fifo_csv_dumper_2045,fifo_intf_2045,cstatus_csv_dumper_2045);
    fifo_csv_dumper_2046 = new("./depth2046.csv");
    cstatus_csv_dumper_2046 = new("./chan_status2046.csv");
    fifo_monitor_2046 = new(fifo_csv_dumper_2046,fifo_intf_2046,cstatus_csv_dumper_2046);
    fifo_csv_dumper_2047 = new("./depth2047.csv");
    cstatus_csv_dumper_2047 = new("./chan_status2047.csv");
    fifo_monitor_2047 = new(fifo_csv_dumper_2047,fifo_intf_2047,cstatus_csv_dumper_2047);
    fifo_csv_dumper_2048 = new("./depth2048.csv");
    cstatus_csv_dumper_2048 = new("./chan_status2048.csv");
    fifo_monitor_2048 = new(fifo_csv_dumper_2048,fifo_intf_2048,cstatus_csv_dumper_2048);
    fifo_csv_dumper_2049 = new("./depth2049.csv");
    cstatus_csv_dumper_2049 = new("./chan_status2049.csv");
    fifo_monitor_2049 = new(fifo_csv_dumper_2049,fifo_intf_2049,cstatus_csv_dumper_2049);
    fifo_csv_dumper_2050 = new("./depth2050.csv");
    cstatus_csv_dumper_2050 = new("./chan_status2050.csv");
    fifo_monitor_2050 = new(fifo_csv_dumper_2050,fifo_intf_2050,cstatus_csv_dumper_2050);
    fifo_csv_dumper_2051 = new("./depth2051.csv");
    cstatus_csv_dumper_2051 = new("./chan_status2051.csv");
    fifo_monitor_2051 = new(fifo_csv_dumper_2051,fifo_intf_2051,cstatus_csv_dumper_2051);
    fifo_csv_dumper_2052 = new("./depth2052.csv");
    cstatus_csv_dumper_2052 = new("./chan_status2052.csv");
    fifo_monitor_2052 = new(fifo_csv_dumper_2052,fifo_intf_2052,cstatus_csv_dumper_2052);
    fifo_csv_dumper_2053 = new("./depth2053.csv");
    cstatus_csv_dumper_2053 = new("./chan_status2053.csv");
    fifo_monitor_2053 = new(fifo_csv_dumper_2053,fifo_intf_2053,cstatus_csv_dumper_2053);
    fifo_csv_dumper_2054 = new("./depth2054.csv");
    cstatus_csv_dumper_2054 = new("./chan_status2054.csv");
    fifo_monitor_2054 = new(fifo_csv_dumper_2054,fifo_intf_2054,cstatus_csv_dumper_2054);
    fifo_csv_dumper_2055 = new("./depth2055.csv");
    cstatus_csv_dumper_2055 = new("./chan_status2055.csv");
    fifo_monitor_2055 = new(fifo_csv_dumper_2055,fifo_intf_2055,cstatus_csv_dumper_2055);
    fifo_csv_dumper_2056 = new("./depth2056.csv");
    cstatus_csv_dumper_2056 = new("./chan_status2056.csv");
    fifo_monitor_2056 = new(fifo_csv_dumper_2056,fifo_intf_2056,cstatus_csv_dumper_2056);
    fifo_csv_dumper_2057 = new("./depth2057.csv");
    cstatus_csv_dumper_2057 = new("./chan_status2057.csv");
    fifo_monitor_2057 = new(fifo_csv_dumper_2057,fifo_intf_2057,cstatus_csv_dumper_2057);
    fifo_csv_dumper_2058 = new("./depth2058.csv");
    cstatus_csv_dumper_2058 = new("./chan_status2058.csv");
    fifo_monitor_2058 = new(fifo_csv_dumper_2058,fifo_intf_2058,cstatus_csv_dumper_2058);
    fifo_csv_dumper_2059 = new("./depth2059.csv");
    cstatus_csv_dumper_2059 = new("./chan_status2059.csv");
    fifo_monitor_2059 = new(fifo_csv_dumper_2059,fifo_intf_2059,cstatus_csv_dumper_2059);
    fifo_csv_dumper_2060 = new("./depth2060.csv");
    cstatus_csv_dumper_2060 = new("./chan_status2060.csv");
    fifo_monitor_2060 = new(fifo_csv_dumper_2060,fifo_intf_2060,cstatus_csv_dumper_2060);
    fifo_csv_dumper_2061 = new("./depth2061.csv");
    cstatus_csv_dumper_2061 = new("./chan_status2061.csv");
    fifo_monitor_2061 = new(fifo_csv_dumper_2061,fifo_intf_2061,cstatus_csv_dumper_2061);
    fifo_csv_dumper_2062 = new("./depth2062.csv");
    cstatus_csv_dumper_2062 = new("./chan_status2062.csv");
    fifo_monitor_2062 = new(fifo_csv_dumper_2062,fifo_intf_2062,cstatus_csv_dumper_2062);
    fifo_csv_dumper_2063 = new("./depth2063.csv");
    cstatus_csv_dumper_2063 = new("./chan_status2063.csv");
    fifo_monitor_2063 = new(fifo_csv_dumper_2063,fifo_intf_2063,cstatus_csv_dumper_2063);
    fifo_csv_dumper_2064 = new("./depth2064.csv");
    cstatus_csv_dumper_2064 = new("./chan_status2064.csv");
    fifo_monitor_2064 = new(fifo_csv_dumper_2064,fifo_intf_2064,cstatus_csv_dumper_2064);
    fifo_csv_dumper_2065 = new("./depth2065.csv");
    cstatus_csv_dumper_2065 = new("./chan_status2065.csv");
    fifo_monitor_2065 = new(fifo_csv_dumper_2065,fifo_intf_2065,cstatus_csv_dumper_2065);
    fifo_csv_dumper_2066 = new("./depth2066.csv");
    cstatus_csv_dumper_2066 = new("./chan_status2066.csv");
    fifo_monitor_2066 = new(fifo_csv_dumper_2066,fifo_intf_2066,cstatus_csv_dumper_2066);
    fifo_csv_dumper_2067 = new("./depth2067.csv");
    cstatus_csv_dumper_2067 = new("./chan_status2067.csv");
    fifo_monitor_2067 = new(fifo_csv_dumper_2067,fifo_intf_2067,cstatus_csv_dumper_2067);
    fifo_csv_dumper_2068 = new("./depth2068.csv");
    cstatus_csv_dumper_2068 = new("./chan_status2068.csv");
    fifo_monitor_2068 = new(fifo_csv_dumper_2068,fifo_intf_2068,cstatus_csv_dumper_2068);
    fifo_csv_dumper_2069 = new("./depth2069.csv");
    cstatus_csv_dumper_2069 = new("./chan_status2069.csv");
    fifo_monitor_2069 = new(fifo_csv_dumper_2069,fifo_intf_2069,cstatus_csv_dumper_2069);
    fifo_csv_dumper_2070 = new("./depth2070.csv");
    cstatus_csv_dumper_2070 = new("./chan_status2070.csv");
    fifo_monitor_2070 = new(fifo_csv_dumper_2070,fifo_intf_2070,cstatus_csv_dumper_2070);
    fifo_csv_dumper_2071 = new("./depth2071.csv");
    cstatus_csv_dumper_2071 = new("./chan_status2071.csv");
    fifo_monitor_2071 = new(fifo_csv_dumper_2071,fifo_intf_2071,cstatus_csv_dumper_2071);
    fifo_csv_dumper_2072 = new("./depth2072.csv");
    cstatus_csv_dumper_2072 = new("./chan_status2072.csv");
    fifo_monitor_2072 = new(fifo_csv_dumper_2072,fifo_intf_2072,cstatus_csv_dumper_2072);
    fifo_csv_dumper_2073 = new("./depth2073.csv");
    cstatus_csv_dumper_2073 = new("./chan_status2073.csv");
    fifo_monitor_2073 = new(fifo_csv_dumper_2073,fifo_intf_2073,cstatus_csv_dumper_2073);
    fifo_csv_dumper_2074 = new("./depth2074.csv");
    cstatus_csv_dumper_2074 = new("./chan_status2074.csv");
    fifo_monitor_2074 = new(fifo_csv_dumper_2074,fifo_intf_2074,cstatus_csv_dumper_2074);
    fifo_csv_dumper_2075 = new("./depth2075.csv");
    cstatus_csv_dumper_2075 = new("./chan_status2075.csv");
    fifo_monitor_2075 = new(fifo_csv_dumper_2075,fifo_intf_2075,cstatus_csv_dumper_2075);
    fifo_csv_dumper_2076 = new("./depth2076.csv");
    cstatus_csv_dumper_2076 = new("./chan_status2076.csv");
    fifo_monitor_2076 = new(fifo_csv_dumper_2076,fifo_intf_2076,cstatus_csv_dumper_2076);
    fifo_csv_dumper_2077 = new("./depth2077.csv");
    cstatus_csv_dumper_2077 = new("./chan_status2077.csv");
    fifo_monitor_2077 = new(fifo_csv_dumper_2077,fifo_intf_2077,cstatus_csv_dumper_2077);
    fifo_csv_dumper_2078 = new("./depth2078.csv");
    cstatus_csv_dumper_2078 = new("./chan_status2078.csv");
    fifo_monitor_2078 = new(fifo_csv_dumper_2078,fifo_intf_2078,cstatus_csv_dumper_2078);
    fifo_csv_dumper_2079 = new("./depth2079.csv");
    cstatus_csv_dumper_2079 = new("./chan_status2079.csv");
    fifo_monitor_2079 = new(fifo_csv_dumper_2079,fifo_intf_2079,cstatus_csv_dumper_2079);
    fifo_csv_dumper_2080 = new("./depth2080.csv");
    cstatus_csv_dumper_2080 = new("./chan_status2080.csv");
    fifo_monitor_2080 = new(fifo_csv_dumper_2080,fifo_intf_2080,cstatus_csv_dumper_2080);
    fifo_csv_dumper_2081 = new("./depth2081.csv");
    cstatus_csv_dumper_2081 = new("./chan_status2081.csv");
    fifo_monitor_2081 = new(fifo_csv_dumper_2081,fifo_intf_2081,cstatus_csv_dumper_2081);
    fifo_csv_dumper_2082 = new("./depth2082.csv");
    cstatus_csv_dumper_2082 = new("./chan_status2082.csv");
    fifo_monitor_2082 = new(fifo_csv_dumper_2082,fifo_intf_2082,cstatus_csv_dumper_2082);
    fifo_csv_dumper_2083 = new("./depth2083.csv");
    cstatus_csv_dumper_2083 = new("./chan_status2083.csv");
    fifo_monitor_2083 = new(fifo_csv_dumper_2083,fifo_intf_2083,cstatus_csv_dumper_2083);
    fifo_csv_dumper_2084 = new("./depth2084.csv");
    cstatus_csv_dumper_2084 = new("./chan_status2084.csv");
    fifo_monitor_2084 = new(fifo_csv_dumper_2084,fifo_intf_2084,cstatus_csv_dumper_2084);
    fifo_csv_dumper_2085 = new("./depth2085.csv");
    cstatus_csv_dumper_2085 = new("./chan_status2085.csv");
    fifo_monitor_2085 = new(fifo_csv_dumper_2085,fifo_intf_2085,cstatus_csv_dumper_2085);
    fifo_csv_dumper_2086 = new("./depth2086.csv");
    cstatus_csv_dumper_2086 = new("./chan_status2086.csv");
    fifo_monitor_2086 = new(fifo_csv_dumper_2086,fifo_intf_2086,cstatus_csv_dumper_2086);
    fifo_csv_dumper_2087 = new("./depth2087.csv");
    cstatus_csv_dumper_2087 = new("./chan_status2087.csv");
    fifo_monitor_2087 = new(fifo_csv_dumper_2087,fifo_intf_2087,cstatus_csv_dumper_2087);
    fifo_csv_dumper_2088 = new("./depth2088.csv");
    cstatus_csv_dumper_2088 = new("./chan_status2088.csv");
    fifo_monitor_2088 = new(fifo_csv_dumper_2088,fifo_intf_2088,cstatus_csv_dumper_2088);
    fifo_csv_dumper_2089 = new("./depth2089.csv");
    cstatus_csv_dumper_2089 = new("./chan_status2089.csv");
    fifo_monitor_2089 = new(fifo_csv_dumper_2089,fifo_intf_2089,cstatus_csv_dumper_2089);
    fifo_csv_dumper_2090 = new("./depth2090.csv");
    cstatus_csv_dumper_2090 = new("./chan_status2090.csv");
    fifo_monitor_2090 = new(fifo_csv_dumper_2090,fifo_intf_2090,cstatus_csv_dumper_2090);
    fifo_csv_dumper_2091 = new("./depth2091.csv");
    cstatus_csv_dumper_2091 = new("./chan_status2091.csv");
    fifo_monitor_2091 = new(fifo_csv_dumper_2091,fifo_intf_2091,cstatus_csv_dumper_2091);
    fifo_csv_dumper_2092 = new("./depth2092.csv");
    cstatus_csv_dumper_2092 = new("./chan_status2092.csv");
    fifo_monitor_2092 = new(fifo_csv_dumper_2092,fifo_intf_2092,cstatus_csv_dumper_2092);
    fifo_csv_dumper_2093 = new("./depth2093.csv");
    cstatus_csv_dumper_2093 = new("./chan_status2093.csv");
    fifo_monitor_2093 = new(fifo_csv_dumper_2093,fifo_intf_2093,cstatus_csv_dumper_2093);
    fifo_csv_dumper_2094 = new("./depth2094.csv");
    cstatus_csv_dumper_2094 = new("./chan_status2094.csv");
    fifo_monitor_2094 = new(fifo_csv_dumper_2094,fifo_intf_2094,cstatus_csv_dumper_2094);
    fifo_csv_dumper_2095 = new("./depth2095.csv");
    cstatus_csv_dumper_2095 = new("./chan_status2095.csv");
    fifo_monitor_2095 = new(fifo_csv_dumper_2095,fifo_intf_2095,cstatus_csv_dumper_2095);
    fifo_csv_dumper_2096 = new("./depth2096.csv");
    cstatus_csv_dumper_2096 = new("./chan_status2096.csv");
    fifo_monitor_2096 = new(fifo_csv_dumper_2096,fifo_intf_2096,cstatus_csv_dumper_2096);
    fifo_csv_dumper_2097 = new("./depth2097.csv");
    cstatus_csv_dumper_2097 = new("./chan_status2097.csv");
    fifo_monitor_2097 = new(fifo_csv_dumper_2097,fifo_intf_2097,cstatus_csv_dumper_2097);
    fifo_csv_dumper_2098 = new("./depth2098.csv");
    cstatus_csv_dumper_2098 = new("./chan_status2098.csv");
    fifo_monitor_2098 = new(fifo_csv_dumper_2098,fifo_intf_2098,cstatus_csv_dumper_2098);
    fifo_csv_dumper_2099 = new("./depth2099.csv");
    cstatus_csv_dumper_2099 = new("./chan_status2099.csv");
    fifo_monitor_2099 = new(fifo_csv_dumper_2099,fifo_intf_2099,cstatus_csv_dumper_2099);
    fifo_csv_dumper_2100 = new("./depth2100.csv");
    cstatus_csv_dumper_2100 = new("./chan_status2100.csv");
    fifo_monitor_2100 = new(fifo_csv_dumper_2100,fifo_intf_2100,cstatus_csv_dumper_2100);
    fifo_csv_dumper_2101 = new("./depth2101.csv");
    cstatus_csv_dumper_2101 = new("./chan_status2101.csv");
    fifo_monitor_2101 = new(fifo_csv_dumper_2101,fifo_intf_2101,cstatus_csv_dumper_2101);
    fifo_csv_dumper_2102 = new("./depth2102.csv");
    cstatus_csv_dumper_2102 = new("./chan_status2102.csv");
    fifo_monitor_2102 = new(fifo_csv_dumper_2102,fifo_intf_2102,cstatus_csv_dumper_2102);
    fifo_csv_dumper_2103 = new("./depth2103.csv");
    cstatus_csv_dumper_2103 = new("./chan_status2103.csv");
    fifo_monitor_2103 = new(fifo_csv_dumper_2103,fifo_intf_2103,cstatus_csv_dumper_2103);
    fifo_csv_dumper_2104 = new("./depth2104.csv");
    cstatus_csv_dumper_2104 = new("./chan_status2104.csv");
    fifo_monitor_2104 = new(fifo_csv_dumper_2104,fifo_intf_2104,cstatus_csv_dumper_2104);
    fifo_csv_dumper_2105 = new("./depth2105.csv");
    cstatus_csv_dumper_2105 = new("./chan_status2105.csv");
    fifo_monitor_2105 = new(fifo_csv_dumper_2105,fifo_intf_2105,cstatus_csv_dumper_2105);
    fifo_csv_dumper_2106 = new("./depth2106.csv");
    cstatus_csv_dumper_2106 = new("./chan_status2106.csv");
    fifo_monitor_2106 = new(fifo_csv_dumper_2106,fifo_intf_2106,cstatus_csv_dumper_2106);
    fifo_csv_dumper_2107 = new("./depth2107.csv");
    cstatus_csv_dumper_2107 = new("./chan_status2107.csv");
    fifo_monitor_2107 = new(fifo_csv_dumper_2107,fifo_intf_2107,cstatus_csv_dumper_2107);
    fifo_csv_dumper_2108 = new("./depth2108.csv");
    cstatus_csv_dumper_2108 = new("./chan_status2108.csv");
    fifo_monitor_2108 = new(fifo_csv_dumper_2108,fifo_intf_2108,cstatus_csv_dumper_2108);
    fifo_csv_dumper_2109 = new("./depth2109.csv");
    cstatus_csv_dumper_2109 = new("./chan_status2109.csv");
    fifo_monitor_2109 = new(fifo_csv_dumper_2109,fifo_intf_2109,cstatus_csv_dumper_2109);
    fifo_csv_dumper_2110 = new("./depth2110.csv");
    cstatus_csv_dumper_2110 = new("./chan_status2110.csv");
    fifo_monitor_2110 = new(fifo_csv_dumper_2110,fifo_intf_2110,cstatus_csv_dumper_2110);
    fifo_csv_dumper_2111 = new("./depth2111.csv");
    cstatus_csv_dumper_2111 = new("./chan_status2111.csv");
    fifo_monitor_2111 = new(fifo_csv_dumper_2111,fifo_intf_2111,cstatus_csv_dumper_2111);
    fifo_csv_dumper_2112 = new("./depth2112.csv");
    cstatus_csv_dumper_2112 = new("./chan_status2112.csv");
    fifo_monitor_2112 = new(fifo_csv_dumper_2112,fifo_intf_2112,cstatus_csv_dumper_2112);
    fifo_csv_dumper_2113 = new("./depth2113.csv");
    cstatus_csv_dumper_2113 = new("./chan_status2113.csv");
    fifo_monitor_2113 = new(fifo_csv_dumper_2113,fifo_intf_2113,cstatus_csv_dumper_2113);
    fifo_csv_dumper_2114 = new("./depth2114.csv");
    cstatus_csv_dumper_2114 = new("./chan_status2114.csv");
    fifo_monitor_2114 = new(fifo_csv_dumper_2114,fifo_intf_2114,cstatus_csv_dumper_2114);
    fifo_csv_dumper_2115 = new("./depth2115.csv");
    cstatus_csv_dumper_2115 = new("./chan_status2115.csv");
    fifo_monitor_2115 = new(fifo_csv_dumper_2115,fifo_intf_2115,cstatus_csv_dumper_2115);
    fifo_csv_dumper_2116 = new("./depth2116.csv");
    cstatus_csv_dumper_2116 = new("./chan_status2116.csv");
    fifo_monitor_2116 = new(fifo_csv_dumper_2116,fifo_intf_2116,cstatus_csv_dumper_2116);
    fifo_csv_dumper_2117 = new("./depth2117.csv");
    cstatus_csv_dumper_2117 = new("./chan_status2117.csv");
    fifo_monitor_2117 = new(fifo_csv_dumper_2117,fifo_intf_2117,cstatus_csv_dumper_2117);
    fifo_csv_dumper_2118 = new("./depth2118.csv");
    cstatus_csv_dumper_2118 = new("./chan_status2118.csv");
    fifo_monitor_2118 = new(fifo_csv_dumper_2118,fifo_intf_2118,cstatus_csv_dumper_2118);
    fifo_csv_dumper_2119 = new("./depth2119.csv");
    cstatus_csv_dumper_2119 = new("./chan_status2119.csv");
    fifo_monitor_2119 = new(fifo_csv_dumper_2119,fifo_intf_2119,cstatus_csv_dumper_2119);
    fifo_csv_dumper_2120 = new("./depth2120.csv");
    cstatus_csv_dumper_2120 = new("./chan_status2120.csv");
    fifo_monitor_2120 = new(fifo_csv_dumper_2120,fifo_intf_2120,cstatus_csv_dumper_2120);
    fifo_csv_dumper_2121 = new("./depth2121.csv");
    cstatus_csv_dumper_2121 = new("./chan_status2121.csv");
    fifo_monitor_2121 = new(fifo_csv_dumper_2121,fifo_intf_2121,cstatus_csv_dumper_2121);
    fifo_csv_dumper_2122 = new("./depth2122.csv");
    cstatus_csv_dumper_2122 = new("./chan_status2122.csv");
    fifo_monitor_2122 = new(fifo_csv_dumper_2122,fifo_intf_2122,cstatus_csv_dumper_2122);
    fifo_csv_dumper_2123 = new("./depth2123.csv");
    cstatus_csv_dumper_2123 = new("./chan_status2123.csv");
    fifo_monitor_2123 = new(fifo_csv_dumper_2123,fifo_intf_2123,cstatus_csv_dumper_2123);
    fifo_csv_dumper_2124 = new("./depth2124.csv");
    cstatus_csv_dumper_2124 = new("./chan_status2124.csv");
    fifo_monitor_2124 = new(fifo_csv_dumper_2124,fifo_intf_2124,cstatus_csv_dumper_2124);
    fifo_csv_dumper_2125 = new("./depth2125.csv");
    cstatus_csv_dumper_2125 = new("./chan_status2125.csv");
    fifo_monitor_2125 = new(fifo_csv_dumper_2125,fifo_intf_2125,cstatus_csv_dumper_2125);
    fifo_csv_dumper_2126 = new("./depth2126.csv");
    cstatus_csv_dumper_2126 = new("./chan_status2126.csv");
    fifo_monitor_2126 = new(fifo_csv_dumper_2126,fifo_intf_2126,cstatus_csv_dumper_2126);
    fifo_csv_dumper_2127 = new("./depth2127.csv");
    cstatus_csv_dumper_2127 = new("./chan_status2127.csv");
    fifo_monitor_2127 = new(fifo_csv_dumper_2127,fifo_intf_2127,cstatus_csv_dumper_2127);
    fifo_csv_dumper_2128 = new("./depth2128.csv");
    cstatus_csv_dumper_2128 = new("./chan_status2128.csv");
    fifo_monitor_2128 = new(fifo_csv_dumper_2128,fifo_intf_2128,cstatus_csv_dumper_2128);
    fifo_csv_dumper_2129 = new("./depth2129.csv");
    cstatus_csv_dumper_2129 = new("./chan_status2129.csv");
    fifo_monitor_2129 = new(fifo_csv_dumper_2129,fifo_intf_2129,cstatus_csv_dumper_2129);
    fifo_csv_dumper_2130 = new("./depth2130.csv");
    cstatus_csv_dumper_2130 = new("./chan_status2130.csv");
    fifo_monitor_2130 = new(fifo_csv_dumper_2130,fifo_intf_2130,cstatus_csv_dumper_2130);
    fifo_csv_dumper_2131 = new("./depth2131.csv");
    cstatus_csv_dumper_2131 = new("./chan_status2131.csv");
    fifo_monitor_2131 = new(fifo_csv_dumper_2131,fifo_intf_2131,cstatus_csv_dumper_2131);
    fifo_csv_dumper_2132 = new("./depth2132.csv");
    cstatus_csv_dumper_2132 = new("./chan_status2132.csv");
    fifo_monitor_2132 = new(fifo_csv_dumper_2132,fifo_intf_2132,cstatus_csv_dumper_2132);
    fifo_csv_dumper_2133 = new("./depth2133.csv");
    cstatus_csv_dumper_2133 = new("./chan_status2133.csv");
    fifo_monitor_2133 = new(fifo_csv_dumper_2133,fifo_intf_2133,cstatus_csv_dumper_2133);
    fifo_csv_dumper_2134 = new("./depth2134.csv");
    cstatus_csv_dumper_2134 = new("./chan_status2134.csv");
    fifo_monitor_2134 = new(fifo_csv_dumper_2134,fifo_intf_2134,cstatus_csv_dumper_2134);
    fifo_csv_dumper_2135 = new("./depth2135.csv");
    cstatus_csv_dumper_2135 = new("./chan_status2135.csv");
    fifo_monitor_2135 = new(fifo_csv_dumper_2135,fifo_intf_2135,cstatus_csv_dumper_2135);
    fifo_csv_dumper_2136 = new("./depth2136.csv");
    cstatus_csv_dumper_2136 = new("./chan_status2136.csv");
    fifo_monitor_2136 = new(fifo_csv_dumper_2136,fifo_intf_2136,cstatus_csv_dumper_2136);
    fifo_csv_dumper_2137 = new("./depth2137.csv");
    cstatus_csv_dumper_2137 = new("./chan_status2137.csv");
    fifo_monitor_2137 = new(fifo_csv_dumper_2137,fifo_intf_2137,cstatus_csv_dumper_2137);
    fifo_csv_dumper_2138 = new("./depth2138.csv");
    cstatus_csv_dumper_2138 = new("./chan_status2138.csv");
    fifo_monitor_2138 = new(fifo_csv_dumper_2138,fifo_intf_2138,cstatus_csv_dumper_2138);
    fifo_csv_dumper_2139 = new("./depth2139.csv");
    cstatus_csv_dumper_2139 = new("./chan_status2139.csv");
    fifo_monitor_2139 = new(fifo_csv_dumper_2139,fifo_intf_2139,cstatus_csv_dumper_2139);
    fifo_csv_dumper_2140 = new("./depth2140.csv");
    cstatus_csv_dumper_2140 = new("./chan_status2140.csv");
    fifo_monitor_2140 = new(fifo_csv_dumper_2140,fifo_intf_2140,cstatus_csv_dumper_2140);
    fifo_csv_dumper_2141 = new("./depth2141.csv");
    cstatus_csv_dumper_2141 = new("./chan_status2141.csv");
    fifo_monitor_2141 = new(fifo_csv_dumper_2141,fifo_intf_2141,cstatus_csv_dumper_2141);
    fifo_csv_dumper_2142 = new("./depth2142.csv");
    cstatus_csv_dumper_2142 = new("./chan_status2142.csv");
    fifo_monitor_2142 = new(fifo_csv_dumper_2142,fifo_intf_2142,cstatus_csv_dumper_2142);
    fifo_csv_dumper_2143 = new("./depth2143.csv");
    cstatus_csv_dumper_2143 = new("./chan_status2143.csv");
    fifo_monitor_2143 = new(fifo_csv_dumper_2143,fifo_intf_2143,cstatus_csv_dumper_2143);
    fifo_csv_dumper_2144 = new("./depth2144.csv");
    cstatus_csv_dumper_2144 = new("./chan_status2144.csv");
    fifo_monitor_2144 = new(fifo_csv_dumper_2144,fifo_intf_2144,cstatus_csv_dumper_2144);
    fifo_csv_dumper_2145 = new("./depth2145.csv");
    cstatus_csv_dumper_2145 = new("./chan_status2145.csv");
    fifo_monitor_2145 = new(fifo_csv_dumper_2145,fifo_intf_2145,cstatus_csv_dumper_2145);
    fifo_csv_dumper_2146 = new("./depth2146.csv");
    cstatus_csv_dumper_2146 = new("./chan_status2146.csv");
    fifo_monitor_2146 = new(fifo_csv_dumper_2146,fifo_intf_2146,cstatus_csv_dumper_2146);
    fifo_csv_dumper_2147 = new("./depth2147.csv");
    cstatus_csv_dumper_2147 = new("./chan_status2147.csv");
    fifo_monitor_2147 = new(fifo_csv_dumper_2147,fifo_intf_2147,cstatus_csv_dumper_2147);
    fifo_csv_dumper_2148 = new("./depth2148.csv");
    cstatus_csv_dumper_2148 = new("./chan_status2148.csv");
    fifo_monitor_2148 = new(fifo_csv_dumper_2148,fifo_intf_2148,cstatus_csv_dumper_2148);
    fifo_csv_dumper_2149 = new("./depth2149.csv");
    cstatus_csv_dumper_2149 = new("./chan_status2149.csv");
    fifo_monitor_2149 = new(fifo_csv_dumper_2149,fifo_intf_2149,cstatus_csv_dumper_2149);
    fifo_csv_dumper_2150 = new("./depth2150.csv");
    cstatus_csv_dumper_2150 = new("./chan_status2150.csv");
    fifo_monitor_2150 = new(fifo_csv_dumper_2150,fifo_intf_2150,cstatus_csv_dumper_2150);
    fifo_csv_dumper_2151 = new("./depth2151.csv");
    cstatus_csv_dumper_2151 = new("./chan_status2151.csv");
    fifo_monitor_2151 = new(fifo_csv_dumper_2151,fifo_intf_2151,cstatus_csv_dumper_2151);
    fifo_csv_dumper_2152 = new("./depth2152.csv");
    cstatus_csv_dumper_2152 = new("./chan_status2152.csv");
    fifo_monitor_2152 = new(fifo_csv_dumper_2152,fifo_intf_2152,cstatus_csv_dumper_2152);
    fifo_csv_dumper_2153 = new("./depth2153.csv");
    cstatus_csv_dumper_2153 = new("./chan_status2153.csv");
    fifo_monitor_2153 = new(fifo_csv_dumper_2153,fifo_intf_2153,cstatus_csv_dumper_2153);
    fifo_csv_dumper_2154 = new("./depth2154.csv");
    cstatus_csv_dumper_2154 = new("./chan_status2154.csv");
    fifo_monitor_2154 = new(fifo_csv_dumper_2154,fifo_intf_2154,cstatus_csv_dumper_2154);
    fifo_csv_dumper_2155 = new("./depth2155.csv");
    cstatus_csv_dumper_2155 = new("./chan_status2155.csv");
    fifo_monitor_2155 = new(fifo_csv_dumper_2155,fifo_intf_2155,cstatus_csv_dumper_2155);
    fifo_csv_dumper_2156 = new("./depth2156.csv");
    cstatus_csv_dumper_2156 = new("./chan_status2156.csv");
    fifo_monitor_2156 = new(fifo_csv_dumper_2156,fifo_intf_2156,cstatus_csv_dumper_2156);
    fifo_csv_dumper_2157 = new("./depth2157.csv");
    cstatus_csv_dumper_2157 = new("./chan_status2157.csv");
    fifo_monitor_2157 = new(fifo_csv_dumper_2157,fifo_intf_2157,cstatus_csv_dumper_2157);
    fifo_csv_dumper_2158 = new("./depth2158.csv");
    cstatus_csv_dumper_2158 = new("./chan_status2158.csv");
    fifo_monitor_2158 = new(fifo_csv_dumper_2158,fifo_intf_2158,cstatus_csv_dumper_2158);
    fifo_csv_dumper_2159 = new("./depth2159.csv");
    cstatus_csv_dumper_2159 = new("./chan_status2159.csv");
    fifo_monitor_2159 = new(fifo_csv_dumper_2159,fifo_intf_2159,cstatus_csv_dumper_2159);
    fifo_csv_dumper_2160 = new("./depth2160.csv");
    cstatus_csv_dumper_2160 = new("./chan_status2160.csv");
    fifo_monitor_2160 = new(fifo_csv_dumper_2160,fifo_intf_2160,cstatus_csv_dumper_2160);
    fifo_csv_dumper_2161 = new("./depth2161.csv");
    cstatus_csv_dumper_2161 = new("./chan_status2161.csv");
    fifo_monitor_2161 = new(fifo_csv_dumper_2161,fifo_intf_2161,cstatus_csv_dumper_2161);
    fifo_csv_dumper_2162 = new("./depth2162.csv");
    cstatus_csv_dumper_2162 = new("./chan_status2162.csv");
    fifo_monitor_2162 = new(fifo_csv_dumper_2162,fifo_intf_2162,cstatus_csv_dumper_2162);
    fifo_csv_dumper_2163 = new("./depth2163.csv");
    cstatus_csv_dumper_2163 = new("./chan_status2163.csv");
    fifo_monitor_2163 = new(fifo_csv_dumper_2163,fifo_intf_2163,cstatus_csv_dumper_2163);
    fifo_csv_dumper_2164 = new("./depth2164.csv");
    cstatus_csv_dumper_2164 = new("./chan_status2164.csv");
    fifo_monitor_2164 = new(fifo_csv_dumper_2164,fifo_intf_2164,cstatus_csv_dumper_2164);
    fifo_csv_dumper_2165 = new("./depth2165.csv");
    cstatus_csv_dumper_2165 = new("./chan_status2165.csv");
    fifo_monitor_2165 = new(fifo_csv_dumper_2165,fifo_intf_2165,cstatus_csv_dumper_2165);
    fifo_csv_dumper_2166 = new("./depth2166.csv");
    cstatus_csv_dumper_2166 = new("./chan_status2166.csv");
    fifo_monitor_2166 = new(fifo_csv_dumper_2166,fifo_intf_2166,cstatus_csv_dumper_2166);
    fifo_csv_dumper_2167 = new("./depth2167.csv");
    cstatus_csv_dumper_2167 = new("./chan_status2167.csv");
    fifo_monitor_2167 = new(fifo_csv_dumper_2167,fifo_intf_2167,cstatus_csv_dumper_2167);
    fifo_csv_dumper_2168 = new("./depth2168.csv");
    cstatus_csv_dumper_2168 = new("./chan_status2168.csv");
    fifo_monitor_2168 = new(fifo_csv_dumper_2168,fifo_intf_2168,cstatus_csv_dumper_2168);
    fifo_csv_dumper_2169 = new("./depth2169.csv");
    cstatus_csv_dumper_2169 = new("./chan_status2169.csv");
    fifo_monitor_2169 = new(fifo_csv_dumper_2169,fifo_intf_2169,cstatus_csv_dumper_2169);
    fifo_csv_dumper_2170 = new("./depth2170.csv");
    cstatus_csv_dumper_2170 = new("./chan_status2170.csv");
    fifo_monitor_2170 = new(fifo_csv_dumper_2170,fifo_intf_2170,cstatus_csv_dumper_2170);
    fifo_csv_dumper_2171 = new("./depth2171.csv");
    cstatus_csv_dumper_2171 = new("./chan_status2171.csv");
    fifo_monitor_2171 = new(fifo_csv_dumper_2171,fifo_intf_2171,cstatus_csv_dumper_2171);
    fifo_csv_dumper_2172 = new("./depth2172.csv");
    cstatus_csv_dumper_2172 = new("./chan_status2172.csv");
    fifo_monitor_2172 = new(fifo_csv_dumper_2172,fifo_intf_2172,cstatus_csv_dumper_2172);
    fifo_csv_dumper_2173 = new("./depth2173.csv");
    cstatus_csv_dumper_2173 = new("./chan_status2173.csv");
    fifo_monitor_2173 = new(fifo_csv_dumper_2173,fifo_intf_2173,cstatus_csv_dumper_2173);
    fifo_csv_dumper_2174 = new("./depth2174.csv");
    cstatus_csv_dumper_2174 = new("./chan_status2174.csv");
    fifo_monitor_2174 = new(fifo_csv_dumper_2174,fifo_intf_2174,cstatus_csv_dumper_2174);
    fifo_csv_dumper_2175 = new("./depth2175.csv");
    cstatus_csv_dumper_2175 = new("./chan_status2175.csv");
    fifo_monitor_2175 = new(fifo_csv_dumper_2175,fifo_intf_2175,cstatus_csv_dumper_2175);
    fifo_csv_dumper_2176 = new("./depth2176.csv");
    cstatus_csv_dumper_2176 = new("./chan_status2176.csv");
    fifo_monitor_2176 = new(fifo_csv_dumper_2176,fifo_intf_2176,cstatus_csv_dumper_2176);
    fifo_csv_dumper_2177 = new("./depth2177.csv");
    cstatus_csv_dumper_2177 = new("./chan_status2177.csv");
    fifo_monitor_2177 = new(fifo_csv_dumper_2177,fifo_intf_2177,cstatus_csv_dumper_2177);
    fifo_csv_dumper_2178 = new("./depth2178.csv");
    cstatus_csv_dumper_2178 = new("./chan_status2178.csv");
    fifo_monitor_2178 = new(fifo_csv_dumper_2178,fifo_intf_2178,cstatus_csv_dumper_2178);
    fifo_csv_dumper_2179 = new("./depth2179.csv");
    cstatus_csv_dumper_2179 = new("./chan_status2179.csv");
    fifo_monitor_2179 = new(fifo_csv_dumper_2179,fifo_intf_2179,cstatus_csv_dumper_2179);
    fifo_csv_dumper_2180 = new("./depth2180.csv");
    cstatus_csv_dumper_2180 = new("./chan_status2180.csv");
    fifo_monitor_2180 = new(fifo_csv_dumper_2180,fifo_intf_2180,cstatus_csv_dumper_2180);
    fifo_csv_dumper_2181 = new("./depth2181.csv");
    cstatus_csv_dumper_2181 = new("./chan_status2181.csv");
    fifo_monitor_2181 = new(fifo_csv_dumper_2181,fifo_intf_2181,cstatus_csv_dumper_2181);
    fifo_csv_dumper_2182 = new("./depth2182.csv");
    cstatus_csv_dumper_2182 = new("./chan_status2182.csv");
    fifo_monitor_2182 = new(fifo_csv_dumper_2182,fifo_intf_2182,cstatus_csv_dumper_2182);
    fifo_csv_dumper_2183 = new("./depth2183.csv");
    cstatus_csv_dumper_2183 = new("./chan_status2183.csv");
    fifo_monitor_2183 = new(fifo_csv_dumper_2183,fifo_intf_2183,cstatus_csv_dumper_2183);
    fifo_csv_dumper_2184 = new("./depth2184.csv");
    cstatus_csv_dumper_2184 = new("./chan_status2184.csv");
    fifo_monitor_2184 = new(fifo_csv_dumper_2184,fifo_intf_2184,cstatus_csv_dumper_2184);
    fifo_csv_dumper_2185 = new("./depth2185.csv");
    cstatus_csv_dumper_2185 = new("./chan_status2185.csv");
    fifo_monitor_2185 = new(fifo_csv_dumper_2185,fifo_intf_2185,cstatus_csv_dumper_2185);
    fifo_csv_dumper_2186 = new("./depth2186.csv");
    cstatus_csv_dumper_2186 = new("./chan_status2186.csv");
    fifo_monitor_2186 = new(fifo_csv_dumper_2186,fifo_intf_2186,cstatus_csv_dumper_2186);
    fifo_csv_dumper_2187 = new("./depth2187.csv");
    cstatus_csv_dumper_2187 = new("./chan_status2187.csv");
    fifo_monitor_2187 = new(fifo_csv_dumper_2187,fifo_intf_2187,cstatus_csv_dumper_2187);
    fifo_csv_dumper_2188 = new("./depth2188.csv");
    cstatus_csv_dumper_2188 = new("./chan_status2188.csv");
    fifo_monitor_2188 = new(fifo_csv_dumper_2188,fifo_intf_2188,cstatus_csv_dumper_2188);
    fifo_csv_dumper_2189 = new("./depth2189.csv");
    cstatus_csv_dumper_2189 = new("./chan_status2189.csv");
    fifo_monitor_2189 = new(fifo_csv_dumper_2189,fifo_intf_2189,cstatus_csv_dumper_2189);
    fifo_csv_dumper_2190 = new("./depth2190.csv");
    cstatus_csv_dumper_2190 = new("./chan_status2190.csv");
    fifo_monitor_2190 = new(fifo_csv_dumper_2190,fifo_intf_2190,cstatus_csv_dumper_2190);
    fifo_csv_dumper_2191 = new("./depth2191.csv");
    cstatus_csv_dumper_2191 = new("./chan_status2191.csv");
    fifo_monitor_2191 = new(fifo_csv_dumper_2191,fifo_intf_2191,cstatus_csv_dumper_2191);
    fifo_csv_dumper_2192 = new("./depth2192.csv");
    cstatus_csv_dumper_2192 = new("./chan_status2192.csv");
    fifo_monitor_2192 = new(fifo_csv_dumper_2192,fifo_intf_2192,cstatus_csv_dumper_2192);
    fifo_csv_dumper_2193 = new("./depth2193.csv");
    cstatus_csv_dumper_2193 = new("./chan_status2193.csv");
    fifo_monitor_2193 = new(fifo_csv_dumper_2193,fifo_intf_2193,cstatus_csv_dumper_2193);
    fifo_csv_dumper_2194 = new("./depth2194.csv");
    cstatus_csv_dumper_2194 = new("./chan_status2194.csv");
    fifo_monitor_2194 = new(fifo_csv_dumper_2194,fifo_intf_2194,cstatus_csv_dumper_2194);
    fifo_csv_dumper_2195 = new("./depth2195.csv");
    cstatus_csv_dumper_2195 = new("./chan_status2195.csv");
    fifo_monitor_2195 = new(fifo_csv_dumper_2195,fifo_intf_2195,cstatus_csv_dumper_2195);
    fifo_csv_dumper_2196 = new("./depth2196.csv");
    cstatus_csv_dumper_2196 = new("./chan_status2196.csv");
    fifo_monitor_2196 = new(fifo_csv_dumper_2196,fifo_intf_2196,cstatus_csv_dumper_2196);
    fifo_csv_dumper_2197 = new("./depth2197.csv");
    cstatus_csv_dumper_2197 = new("./chan_status2197.csv");
    fifo_monitor_2197 = new(fifo_csv_dumper_2197,fifo_intf_2197,cstatus_csv_dumper_2197);
    fifo_csv_dumper_2198 = new("./depth2198.csv");
    cstatus_csv_dumper_2198 = new("./chan_status2198.csv");
    fifo_monitor_2198 = new(fifo_csv_dumper_2198,fifo_intf_2198,cstatus_csv_dumper_2198);
    fifo_csv_dumper_2199 = new("./depth2199.csv");
    cstatus_csv_dumper_2199 = new("./chan_status2199.csv");
    fifo_monitor_2199 = new(fifo_csv_dumper_2199,fifo_intf_2199,cstatus_csv_dumper_2199);
    fifo_csv_dumper_2200 = new("./depth2200.csv");
    cstatus_csv_dumper_2200 = new("./chan_status2200.csv");
    fifo_monitor_2200 = new(fifo_csv_dumper_2200,fifo_intf_2200,cstatus_csv_dumper_2200);
    fifo_csv_dumper_2201 = new("./depth2201.csv");
    cstatus_csv_dumper_2201 = new("./chan_status2201.csv");
    fifo_monitor_2201 = new(fifo_csv_dumper_2201,fifo_intf_2201,cstatus_csv_dumper_2201);
    fifo_csv_dumper_2202 = new("./depth2202.csv");
    cstatus_csv_dumper_2202 = new("./chan_status2202.csv");
    fifo_monitor_2202 = new(fifo_csv_dumper_2202,fifo_intf_2202,cstatus_csv_dumper_2202);
    fifo_csv_dumper_2203 = new("./depth2203.csv");
    cstatus_csv_dumper_2203 = new("./chan_status2203.csv");
    fifo_monitor_2203 = new(fifo_csv_dumper_2203,fifo_intf_2203,cstatus_csv_dumper_2203);
    fifo_csv_dumper_2204 = new("./depth2204.csv");
    cstatus_csv_dumper_2204 = new("./chan_status2204.csv");
    fifo_monitor_2204 = new(fifo_csv_dumper_2204,fifo_intf_2204,cstatus_csv_dumper_2204);
    fifo_csv_dumper_2205 = new("./depth2205.csv");
    cstatus_csv_dumper_2205 = new("./chan_status2205.csv");
    fifo_monitor_2205 = new(fifo_csv_dumper_2205,fifo_intf_2205,cstatus_csv_dumper_2205);
    fifo_csv_dumper_2206 = new("./depth2206.csv");
    cstatus_csv_dumper_2206 = new("./chan_status2206.csv");
    fifo_monitor_2206 = new(fifo_csv_dumper_2206,fifo_intf_2206,cstatus_csv_dumper_2206);
    fifo_csv_dumper_2207 = new("./depth2207.csv");
    cstatus_csv_dumper_2207 = new("./chan_status2207.csv");
    fifo_monitor_2207 = new(fifo_csv_dumper_2207,fifo_intf_2207,cstatus_csv_dumper_2207);
    fifo_csv_dumper_2208 = new("./depth2208.csv");
    cstatus_csv_dumper_2208 = new("./chan_status2208.csv");
    fifo_monitor_2208 = new(fifo_csv_dumper_2208,fifo_intf_2208,cstatus_csv_dumper_2208);
    fifo_csv_dumper_2209 = new("./depth2209.csv");
    cstatus_csv_dumper_2209 = new("./chan_status2209.csv");
    fifo_monitor_2209 = new(fifo_csv_dumper_2209,fifo_intf_2209,cstatus_csv_dumper_2209);
    fifo_csv_dumper_2210 = new("./depth2210.csv");
    cstatus_csv_dumper_2210 = new("./chan_status2210.csv");
    fifo_monitor_2210 = new(fifo_csv_dumper_2210,fifo_intf_2210,cstatus_csv_dumper_2210);
    fifo_csv_dumper_2211 = new("./depth2211.csv");
    cstatus_csv_dumper_2211 = new("./chan_status2211.csv");
    fifo_monitor_2211 = new(fifo_csv_dumper_2211,fifo_intf_2211,cstatus_csv_dumper_2211);
    fifo_csv_dumper_2212 = new("./depth2212.csv");
    cstatus_csv_dumper_2212 = new("./chan_status2212.csv");
    fifo_monitor_2212 = new(fifo_csv_dumper_2212,fifo_intf_2212,cstatus_csv_dumper_2212);
    fifo_csv_dumper_2213 = new("./depth2213.csv");
    cstatus_csv_dumper_2213 = new("./chan_status2213.csv");
    fifo_monitor_2213 = new(fifo_csv_dumper_2213,fifo_intf_2213,cstatus_csv_dumper_2213);
    fifo_csv_dumper_2214 = new("./depth2214.csv");
    cstatus_csv_dumper_2214 = new("./chan_status2214.csv");
    fifo_monitor_2214 = new(fifo_csv_dumper_2214,fifo_intf_2214,cstatus_csv_dumper_2214);
    fifo_csv_dumper_2215 = new("./depth2215.csv");
    cstatus_csv_dumper_2215 = new("./chan_status2215.csv");
    fifo_monitor_2215 = new(fifo_csv_dumper_2215,fifo_intf_2215,cstatus_csv_dumper_2215);
    fifo_csv_dumper_2216 = new("./depth2216.csv");
    cstatus_csv_dumper_2216 = new("./chan_status2216.csv");
    fifo_monitor_2216 = new(fifo_csv_dumper_2216,fifo_intf_2216,cstatus_csv_dumper_2216);
    fifo_csv_dumper_2217 = new("./depth2217.csv");
    cstatus_csv_dumper_2217 = new("./chan_status2217.csv");
    fifo_monitor_2217 = new(fifo_csv_dumper_2217,fifo_intf_2217,cstatus_csv_dumper_2217);
    fifo_csv_dumper_2218 = new("./depth2218.csv");
    cstatus_csv_dumper_2218 = new("./chan_status2218.csv");
    fifo_monitor_2218 = new(fifo_csv_dumper_2218,fifo_intf_2218,cstatus_csv_dumper_2218);
    fifo_csv_dumper_2219 = new("./depth2219.csv");
    cstatus_csv_dumper_2219 = new("./chan_status2219.csv");
    fifo_monitor_2219 = new(fifo_csv_dumper_2219,fifo_intf_2219,cstatus_csv_dumper_2219);
    fifo_csv_dumper_2220 = new("./depth2220.csv");
    cstatus_csv_dumper_2220 = new("./chan_status2220.csv");
    fifo_monitor_2220 = new(fifo_csv_dumper_2220,fifo_intf_2220,cstatus_csv_dumper_2220);
    fifo_csv_dumper_2221 = new("./depth2221.csv");
    cstatus_csv_dumper_2221 = new("./chan_status2221.csv");
    fifo_monitor_2221 = new(fifo_csv_dumper_2221,fifo_intf_2221,cstatus_csv_dumper_2221);
    fifo_csv_dumper_2222 = new("./depth2222.csv");
    cstatus_csv_dumper_2222 = new("./chan_status2222.csv");
    fifo_monitor_2222 = new(fifo_csv_dumper_2222,fifo_intf_2222,cstatus_csv_dumper_2222);
    fifo_csv_dumper_2223 = new("./depth2223.csv");
    cstatus_csv_dumper_2223 = new("./chan_status2223.csv");
    fifo_monitor_2223 = new(fifo_csv_dumper_2223,fifo_intf_2223,cstatus_csv_dumper_2223);
    fifo_csv_dumper_2224 = new("./depth2224.csv");
    cstatus_csv_dumper_2224 = new("./chan_status2224.csv");
    fifo_monitor_2224 = new(fifo_csv_dumper_2224,fifo_intf_2224,cstatus_csv_dumper_2224);
    fifo_csv_dumper_2225 = new("./depth2225.csv");
    cstatus_csv_dumper_2225 = new("./chan_status2225.csv");
    fifo_monitor_2225 = new(fifo_csv_dumper_2225,fifo_intf_2225,cstatus_csv_dumper_2225);
    fifo_csv_dumper_2226 = new("./depth2226.csv");
    cstatus_csv_dumper_2226 = new("./chan_status2226.csv");
    fifo_monitor_2226 = new(fifo_csv_dumper_2226,fifo_intf_2226,cstatus_csv_dumper_2226);
    fifo_csv_dumper_2227 = new("./depth2227.csv");
    cstatus_csv_dumper_2227 = new("./chan_status2227.csv");
    fifo_monitor_2227 = new(fifo_csv_dumper_2227,fifo_intf_2227,cstatus_csv_dumper_2227);
    fifo_csv_dumper_2228 = new("./depth2228.csv");
    cstatus_csv_dumper_2228 = new("./chan_status2228.csv");
    fifo_monitor_2228 = new(fifo_csv_dumper_2228,fifo_intf_2228,cstatus_csv_dumper_2228);
    fifo_csv_dumper_2229 = new("./depth2229.csv");
    cstatus_csv_dumper_2229 = new("./chan_status2229.csv");
    fifo_monitor_2229 = new(fifo_csv_dumper_2229,fifo_intf_2229,cstatus_csv_dumper_2229);
    fifo_csv_dumper_2230 = new("./depth2230.csv");
    cstatus_csv_dumper_2230 = new("./chan_status2230.csv");
    fifo_monitor_2230 = new(fifo_csv_dumper_2230,fifo_intf_2230,cstatus_csv_dumper_2230);
    fifo_csv_dumper_2231 = new("./depth2231.csv");
    cstatus_csv_dumper_2231 = new("./chan_status2231.csv");
    fifo_monitor_2231 = new(fifo_csv_dumper_2231,fifo_intf_2231,cstatus_csv_dumper_2231);
    fifo_csv_dumper_2232 = new("./depth2232.csv");
    cstatus_csv_dumper_2232 = new("./chan_status2232.csv");
    fifo_monitor_2232 = new(fifo_csv_dumper_2232,fifo_intf_2232,cstatus_csv_dumper_2232);
    fifo_csv_dumper_2233 = new("./depth2233.csv");
    cstatus_csv_dumper_2233 = new("./chan_status2233.csv");
    fifo_monitor_2233 = new(fifo_csv_dumper_2233,fifo_intf_2233,cstatus_csv_dumper_2233);
    fifo_csv_dumper_2234 = new("./depth2234.csv");
    cstatus_csv_dumper_2234 = new("./chan_status2234.csv");
    fifo_monitor_2234 = new(fifo_csv_dumper_2234,fifo_intf_2234,cstatus_csv_dumper_2234);
    fifo_csv_dumper_2235 = new("./depth2235.csv");
    cstatus_csv_dumper_2235 = new("./chan_status2235.csv");
    fifo_monitor_2235 = new(fifo_csv_dumper_2235,fifo_intf_2235,cstatus_csv_dumper_2235);
    fifo_csv_dumper_2236 = new("./depth2236.csv");
    cstatus_csv_dumper_2236 = new("./chan_status2236.csv");
    fifo_monitor_2236 = new(fifo_csv_dumper_2236,fifo_intf_2236,cstatus_csv_dumper_2236);
    fifo_csv_dumper_2237 = new("./depth2237.csv");
    cstatus_csv_dumper_2237 = new("./chan_status2237.csv");
    fifo_monitor_2237 = new(fifo_csv_dumper_2237,fifo_intf_2237,cstatus_csv_dumper_2237);
    fifo_csv_dumper_2238 = new("./depth2238.csv");
    cstatus_csv_dumper_2238 = new("./chan_status2238.csv");
    fifo_monitor_2238 = new(fifo_csv_dumper_2238,fifo_intf_2238,cstatus_csv_dumper_2238);
    fifo_csv_dumper_2239 = new("./depth2239.csv");
    cstatus_csv_dumper_2239 = new("./chan_status2239.csv");
    fifo_monitor_2239 = new(fifo_csv_dumper_2239,fifo_intf_2239,cstatus_csv_dumper_2239);
    fifo_csv_dumper_2240 = new("./depth2240.csv");
    cstatus_csv_dumper_2240 = new("./chan_status2240.csv");
    fifo_monitor_2240 = new(fifo_csv_dumper_2240,fifo_intf_2240,cstatus_csv_dumper_2240);
    fifo_csv_dumper_2241 = new("./depth2241.csv");
    cstatus_csv_dumper_2241 = new("./chan_status2241.csv");
    fifo_monitor_2241 = new(fifo_csv_dumper_2241,fifo_intf_2241,cstatus_csv_dumper_2241);
    fifo_csv_dumper_2242 = new("./depth2242.csv");
    cstatus_csv_dumper_2242 = new("./chan_status2242.csv");
    fifo_monitor_2242 = new(fifo_csv_dumper_2242,fifo_intf_2242,cstatus_csv_dumper_2242);
    fifo_csv_dumper_2243 = new("./depth2243.csv");
    cstatus_csv_dumper_2243 = new("./chan_status2243.csv");
    fifo_monitor_2243 = new(fifo_csv_dumper_2243,fifo_intf_2243,cstatus_csv_dumper_2243);
    fifo_csv_dumper_2244 = new("./depth2244.csv");
    cstatus_csv_dumper_2244 = new("./chan_status2244.csv");
    fifo_monitor_2244 = new(fifo_csv_dumper_2244,fifo_intf_2244,cstatus_csv_dumper_2244);
    fifo_csv_dumper_2245 = new("./depth2245.csv");
    cstatus_csv_dumper_2245 = new("./chan_status2245.csv");
    fifo_monitor_2245 = new(fifo_csv_dumper_2245,fifo_intf_2245,cstatus_csv_dumper_2245);
    fifo_csv_dumper_2246 = new("./depth2246.csv");
    cstatus_csv_dumper_2246 = new("./chan_status2246.csv");
    fifo_monitor_2246 = new(fifo_csv_dumper_2246,fifo_intf_2246,cstatus_csv_dumper_2246);
    fifo_csv_dumper_2247 = new("./depth2247.csv");
    cstatus_csv_dumper_2247 = new("./chan_status2247.csv");
    fifo_monitor_2247 = new(fifo_csv_dumper_2247,fifo_intf_2247,cstatus_csv_dumper_2247);
    fifo_csv_dumper_2248 = new("./depth2248.csv");
    cstatus_csv_dumper_2248 = new("./chan_status2248.csv");
    fifo_monitor_2248 = new(fifo_csv_dumper_2248,fifo_intf_2248,cstatus_csv_dumper_2248);
    fifo_csv_dumper_2249 = new("./depth2249.csv");
    cstatus_csv_dumper_2249 = new("./chan_status2249.csv");
    fifo_monitor_2249 = new(fifo_csv_dumper_2249,fifo_intf_2249,cstatus_csv_dumper_2249);
    fifo_csv_dumper_2250 = new("./depth2250.csv");
    cstatus_csv_dumper_2250 = new("./chan_status2250.csv");
    fifo_monitor_2250 = new(fifo_csv_dumper_2250,fifo_intf_2250,cstatus_csv_dumper_2250);
    fifo_csv_dumper_2251 = new("./depth2251.csv");
    cstatus_csv_dumper_2251 = new("./chan_status2251.csv");
    fifo_monitor_2251 = new(fifo_csv_dumper_2251,fifo_intf_2251,cstatus_csv_dumper_2251);
    fifo_csv_dumper_2252 = new("./depth2252.csv");
    cstatus_csv_dumper_2252 = new("./chan_status2252.csv");
    fifo_monitor_2252 = new(fifo_csv_dumper_2252,fifo_intf_2252,cstatus_csv_dumper_2252);
    fifo_csv_dumper_2253 = new("./depth2253.csv");
    cstatus_csv_dumper_2253 = new("./chan_status2253.csv");
    fifo_monitor_2253 = new(fifo_csv_dumper_2253,fifo_intf_2253,cstatus_csv_dumper_2253);
    fifo_csv_dumper_2254 = new("./depth2254.csv");
    cstatus_csv_dumper_2254 = new("./chan_status2254.csv");
    fifo_monitor_2254 = new(fifo_csv_dumper_2254,fifo_intf_2254,cstatus_csv_dumper_2254);
    fifo_csv_dumper_2255 = new("./depth2255.csv");
    cstatus_csv_dumper_2255 = new("./chan_status2255.csv");
    fifo_monitor_2255 = new(fifo_csv_dumper_2255,fifo_intf_2255,cstatus_csv_dumper_2255);
    fifo_csv_dumper_2256 = new("./depth2256.csv");
    cstatus_csv_dumper_2256 = new("./chan_status2256.csv");
    fifo_monitor_2256 = new(fifo_csv_dumper_2256,fifo_intf_2256,cstatus_csv_dumper_2256);
    fifo_csv_dumper_2257 = new("./depth2257.csv");
    cstatus_csv_dumper_2257 = new("./chan_status2257.csv");
    fifo_monitor_2257 = new(fifo_csv_dumper_2257,fifo_intf_2257,cstatus_csv_dumper_2257);
    fifo_csv_dumper_2258 = new("./depth2258.csv");
    cstatus_csv_dumper_2258 = new("./chan_status2258.csv");
    fifo_monitor_2258 = new(fifo_csv_dumper_2258,fifo_intf_2258,cstatus_csv_dumper_2258);
    fifo_csv_dumper_2259 = new("./depth2259.csv");
    cstatus_csv_dumper_2259 = new("./chan_status2259.csv");
    fifo_monitor_2259 = new(fifo_csv_dumper_2259,fifo_intf_2259,cstatus_csv_dumper_2259);
    fifo_csv_dumper_2260 = new("./depth2260.csv");
    cstatus_csv_dumper_2260 = new("./chan_status2260.csv");
    fifo_monitor_2260 = new(fifo_csv_dumper_2260,fifo_intf_2260,cstatus_csv_dumper_2260);
    fifo_csv_dumper_2261 = new("./depth2261.csv");
    cstatus_csv_dumper_2261 = new("./chan_status2261.csv");
    fifo_monitor_2261 = new(fifo_csv_dumper_2261,fifo_intf_2261,cstatus_csv_dumper_2261);
    fifo_csv_dumper_2262 = new("./depth2262.csv");
    cstatus_csv_dumper_2262 = new("./chan_status2262.csv");
    fifo_monitor_2262 = new(fifo_csv_dumper_2262,fifo_intf_2262,cstatus_csv_dumper_2262);
    fifo_csv_dumper_2263 = new("./depth2263.csv");
    cstatus_csv_dumper_2263 = new("./chan_status2263.csv");
    fifo_monitor_2263 = new(fifo_csv_dumper_2263,fifo_intf_2263,cstatus_csv_dumper_2263);
    fifo_csv_dumper_2264 = new("./depth2264.csv");
    cstatus_csv_dumper_2264 = new("./chan_status2264.csv");
    fifo_monitor_2264 = new(fifo_csv_dumper_2264,fifo_intf_2264,cstatus_csv_dumper_2264);
    fifo_csv_dumper_2265 = new("./depth2265.csv");
    cstatus_csv_dumper_2265 = new("./chan_status2265.csv");
    fifo_monitor_2265 = new(fifo_csv_dumper_2265,fifo_intf_2265,cstatus_csv_dumper_2265);
    fifo_csv_dumper_2266 = new("./depth2266.csv");
    cstatus_csv_dumper_2266 = new("./chan_status2266.csv");
    fifo_monitor_2266 = new(fifo_csv_dumper_2266,fifo_intf_2266,cstatus_csv_dumper_2266);
    fifo_csv_dumper_2267 = new("./depth2267.csv");
    cstatus_csv_dumper_2267 = new("./chan_status2267.csv");
    fifo_monitor_2267 = new(fifo_csv_dumper_2267,fifo_intf_2267,cstatus_csv_dumper_2267);
    fifo_csv_dumper_2268 = new("./depth2268.csv");
    cstatus_csv_dumper_2268 = new("./chan_status2268.csv");
    fifo_monitor_2268 = new(fifo_csv_dumper_2268,fifo_intf_2268,cstatus_csv_dumper_2268);
    fifo_csv_dumper_2269 = new("./depth2269.csv");
    cstatus_csv_dumper_2269 = new("./chan_status2269.csv");
    fifo_monitor_2269 = new(fifo_csv_dumper_2269,fifo_intf_2269,cstatus_csv_dumper_2269);
    fifo_csv_dumper_2270 = new("./depth2270.csv");
    cstatus_csv_dumper_2270 = new("./chan_status2270.csv");
    fifo_monitor_2270 = new(fifo_csv_dumper_2270,fifo_intf_2270,cstatus_csv_dumper_2270);
    fifo_csv_dumper_2271 = new("./depth2271.csv");
    cstatus_csv_dumper_2271 = new("./chan_status2271.csv");
    fifo_monitor_2271 = new(fifo_csv_dumper_2271,fifo_intf_2271,cstatus_csv_dumper_2271);
    fifo_csv_dumper_2272 = new("./depth2272.csv");
    cstatus_csv_dumper_2272 = new("./chan_status2272.csv");
    fifo_monitor_2272 = new(fifo_csv_dumper_2272,fifo_intf_2272,cstatus_csv_dumper_2272);
    fifo_csv_dumper_2273 = new("./depth2273.csv");
    cstatus_csv_dumper_2273 = new("./chan_status2273.csv");
    fifo_monitor_2273 = new(fifo_csv_dumper_2273,fifo_intf_2273,cstatus_csv_dumper_2273);
    fifo_csv_dumper_2274 = new("./depth2274.csv");
    cstatus_csv_dumper_2274 = new("./chan_status2274.csv");
    fifo_monitor_2274 = new(fifo_csv_dumper_2274,fifo_intf_2274,cstatus_csv_dumper_2274);
    fifo_csv_dumper_2275 = new("./depth2275.csv");
    cstatus_csv_dumper_2275 = new("./chan_status2275.csv");
    fifo_monitor_2275 = new(fifo_csv_dumper_2275,fifo_intf_2275,cstatus_csv_dumper_2275);
    fifo_csv_dumper_2276 = new("./depth2276.csv");
    cstatus_csv_dumper_2276 = new("./chan_status2276.csv");
    fifo_monitor_2276 = new(fifo_csv_dumper_2276,fifo_intf_2276,cstatus_csv_dumper_2276);
    fifo_csv_dumper_2277 = new("./depth2277.csv");
    cstatus_csv_dumper_2277 = new("./chan_status2277.csv");
    fifo_monitor_2277 = new(fifo_csv_dumper_2277,fifo_intf_2277,cstatus_csv_dumper_2277);
    fifo_csv_dumper_2278 = new("./depth2278.csv");
    cstatus_csv_dumper_2278 = new("./chan_status2278.csv");
    fifo_monitor_2278 = new(fifo_csv_dumper_2278,fifo_intf_2278,cstatus_csv_dumper_2278);
    fifo_csv_dumper_2279 = new("./depth2279.csv");
    cstatus_csv_dumper_2279 = new("./chan_status2279.csv");
    fifo_monitor_2279 = new(fifo_csv_dumper_2279,fifo_intf_2279,cstatus_csv_dumper_2279);
    fifo_csv_dumper_2280 = new("./depth2280.csv");
    cstatus_csv_dumper_2280 = new("./chan_status2280.csv");
    fifo_monitor_2280 = new(fifo_csv_dumper_2280,fifo_intf_2280,cstatus_csv_dumper_2280);
    fifo_csv_dumper_2281 = new("./depth2281.csv");
    cstatus_csv_dumper_2281 = new("./chan_status2281.csv");
    fifo_monitor_2281 = new(fifo_csv_dumper_2281,fifo_intf_2281,cstatus_csv_dumper_2281);
    fifo_csv_dumper_2282 = new("./depth2282.csv");
    cstatus_csv_dumper_2282 = new("./chan_status2282.csv");
    fifo_monitor_2282 = new(fifo_csv_dumper_2282,fifo_intf_2282,cstatus_csv_dumper_2282);
    fifo_csv_dumper_2283 = new("./depth2283.csv");
    cstatus_csv_dumper_2283 = new("./chan_status2283.csv");
    fifo_monitor_2283 = new(fifo_csv_dumper_2283,fifo_intf_2283,cstatus_csv_dumper_2283);
    fifo_csv_dumper_2284 = new("./depth2284.csv");
    cstatus_csv_dumper_2284 = new("./chan_status2284.csv");
    fifo_monitor_2284 = new(fifo_csv_dumper_2284,fifo_intf_2284,cstatus_csv_dumper_2284);
    fifo_csv_dumper_2285 = new("./depth2285.csv");
    cstatus_csv_dumper_2285 = new("./chan_status2285.csv");
    fifo_monitor_2285 = new(fifo_csv_dumper_2285,fifo_intf_2285,cstatus_csv_dumper_2285);
    fifo_csv_dumper_2286 = new("./depth2286.csv");
    cstatus_csv_dumper_2286 = new("./chan_status2286.csv");
    fifo_monitor_2286 = new(fifo_csv_dumper_2286,fifo_intf_2286,cstatus_csv_dumper_2286);
    fifo_csv_dumper_2287 = new("./depth2287.csv");
    cstatus_csv_dumper_2287 = new("./chan_status2287.csv");
    fifo_monitor_2287 = new(fifo_csv_dumper_2287,fifo_intf_2287,cstatus_csv_dumper_2287);
    fifo_csv_dumper_2288 = new("./depth2288.csv");
    cstatus_csv_dumper_2288 = new("./chan_status2288.csv");
    fifo_monitor_2288 = new(fifo_csv_dumper_2288,fifo_intf_2288,cstatus_csv_dumper_2288);
    fifo_csv_dumper_2289 = new("./depth2289.csv");
    cstatus_csv_dumper_2289 = new("./chan_status2289.csv");
    fifo_monitor_2289 = new(fifo_csv_dumper_2289,fifo_intf_2289,cstatus_csv_dumper_2289);
    fifo_csv_dumper_2290 = new("./depth2290.csv");
    cstatus_csv_dumper_2290 = new("./chan_status2290.csv");
    fifo_monitor_2290 = new(fifo_csv_dumper_2290,fifo_intf_2290,cstatus_csv_dumper_2290);
    fifo_csv_dumper_2291 = new("./depth2291.csv");
    cstatus_csv_dumper_2291 = new("./chan_status2291.csv");
    fifo_monitor_2291 = new(fifo_csv_dumper_2291,fifo_intf_2291,cstatus_csv_dumper_2291);
    fifo_csv_dumper_2292 = new("./depth2292.csv");
    cstatus_csv_dumper_2292 = new("./chan_status2292.csv");
    fifo_monitor_2292 = new(fifo_csv_dumper_2292,fifo_intf_2292,cstatus_csv_dumper_2292);
    fifo_csv_dumper_2293 = new("./depth2293.csv");
    cstatus_csv_dumper_2293 = new("./chan_status2293.csv");
    fifo_monitor_2293 = new(fifo_csv_dumper_2293,fifo_intf_2293,cstatus_csv_dumper_2293);
    fifo_csv_dumper_2294 = new("./depth2294.csv");
    cstatus_csv_dumper_2294 = new("./chan_status2294.csv");
    fifo_monitor_2294 = new(fifo_csv_dumper_2294,fifo_intf_2294,cstatus_csv_dumper_2294);
    fifo_csv_dumper_2295 = new("./depth2295.csv");
    cstatus_csv_dumper_2295 = new("./chan_status2295.csv");
    fifo_monitor_2295 = new(fifo_csv_dumper_2295,fifo_intf_2295,cstatus_csv_dumper_2295);
    fifo_csv_dumper_2296 = new("./depth2296.csv");
    cstatus_csv_dumper_2296 = new("./chan_status2296.csv");
    fifo_monitor_2296 = new(fifo_csv_dumper_2296,fifo_intf_2296,cstatus_csv_dumper_2296);
    fifo_csv_dumper_2297 = new("./depth2297.csv");
    cstatus_csv_dumper_2297 = new("./chan_status2297.csv");
    fifo_monitor_2297 = new(fifo_csv_dumper_2297,fifo_intf_2297,cstatus_csv_dumper_2297);
    fifo_csv_dumper_2298 = new("./depth2298.csv");
    cstatus_csv_dumper_2298 = new("./chan_status2298.csv");
    fifo_monitor_2298 = new(fifo_csv_dumper_2298,fifo_intf_2298,cstatus_csv_dumper_2298);
    fifo_csv_dumper_2299 = new("./depth2299.csv");
    cstatus_csv_dumper_2299 = new("./chan_status2299.csv");
    fifo_monitor_2299 = new(fifo_csv_dumper_2299,fifo_intf_2299,cstatus_csv_dumper_2299);
    fifo_csv_dumper_2300 = new("./depth2300.csv");
    cstatus_csv_dumper_2300 = new("./chan_status2300.csv");
    fifo_monitor_2300 = new(fifo_csv_dumper_2300,fifo_intf_2300,cstatus_csv_dumper_2300);
    fifo_csv_dumper_2301 = new("./depth2301.csv");
    cstatus_csv_dumper_2301 = new("./chan_status2301.csv");
    fifo_monitor_2301 = new(fifo_csv_dumper_2301,fifo_intf_2301,cstatus_csv_dumper_2301);
    fifo_csv_dumper_2302 = new("./depth2302.csv");
    cstatus_csv_dumper_2302 = new("./chan_status2302.csv");
    fifo_monitor_2302 = new(fifo_csv_dumper_2302,fifo_intf_2302,cstatus_csv_dumper_2302);
    fifo_csv_dumper_2303 = new("./depth2303.csv");
    cstatus_csv_dumper_2303 = new("./chan_status2303.csv");
    fifo_monitor_2303 = new(fifo_csv_dumper_2303,fifo_intf_2303,cstatus_csv_dumper_2303);
    fifo_csv_dumper_2304 = new("./depth2304.csv");
    cstatus_csv_dumper_2304 = new("./chan_status2304.csv");
    fifo_monitor_2304 = new(fifo_csv_dumper_2304,fifo_intf_2304,cstatus_csv_dumper_2304);
    fifo_csv_dumper_2305 = new("./depth2305.csv");
    cstatus_csv_dumper_2305 = new("./chan_status2305.csv");
    fifo_monitor_2305 = new(fifo_csv_dumper_2305,fifo_intf_2305,cstatus_csv_dumper_2305);
    fifo_csv_dumper_2306 = new("./depth2306.csv");
    cstatus_csv_dumper_2306 = new("./chan_status2306.csv");
    fifo_monitor_2306 = new(fifo_csv_dumper_2306,fifo_intf_2306,cstatus_csv_dumper_2306);
    fifo_csv_dumper_2307 = new("./depth2307.csv");
    cstatus_csv_dumper_2307 = new("./chan_status2307.csv");
    fifo_monitor_2307 = new(fifo_csv_dumper_2307,fifo_intf_2307,cstatus_csv_dumper_2307);
    fifo_csv_dumper_2308 = new("./depth2308.csv");
    cstatus_csv_dumper_2308 = new("./chan_status2308.csv");
    fifo_monitor_2308 = new(fifo_csv_dumper_2308,fifo_intf_2308,cstatus_csv_dumper_2308);
    fifo_csv_dumper_2309 = new("./depth2309.csv");
    cstatus_csv_dumper_2309 = new("./chan_status2309.csv");
    fifo_monitor_2309 = new(fifo_csv_dumper_2309,fifo_intf_2309,cstatus_csv_dumper_2309);
    fifo_csv_dumper_2310 = new("./depth2310.csv");
    cstatus_csv_dumper_2310 = new("./chan_status2310.csv");
    fifo_monitor_2310 = new(fifo_csv_dumper_2310,fifo_intf_2310,cstatus_csv_dumper_2310);
    fifo_csv_dumper_2311 = new("./depth2311.csv");
    cstatus_csv_dumper_2311 = new("./chan_status2311.csv");
    fifo_monitor_2311 = new(fifo_csv_dumper_2311,fifo_intf_2311,cstatus_csv_dumper_2311);
    fifo_csv_dumper_2312 = new("./depth2312.csv");
    cstatus_csv_dumper_2312 = new("./chan_status2312.csv");
    fifo_monitor_2312 = new(fifo_csv_dumper_2312,fifo_intf_2312,cstatus_csv_dumper_2312);
    fifo_csv_dumper_2313 = new("./depth2313.csv");
    cstatus_csv_dumper_2313 = new("./chan_status2313.csv");
    fifo_monitor_2313 = new(fifo_csv_dumper_2313,fifo_intf_2313,cstatus_csv_dumper_2313);
    fifo_csv_dumper_2314 = new("./depth2314.csv");
    cstatus_csv_dumper_2314 = new("./chan_status2314.csv");
    fifo_monitor_2314 = new(fifo_csv_dumper_2314,fifo_intf_2314,cstatus_csv_dumper_2314);
    fifo_csv_dumper_2315 = new("./depth2315.csv");
    cstatus_csv_dumper_2315 = new("./chan_status2315.csv");
    fifo_monitor_2315 = new(fifo_csv_dumper_2315,fifo_intf_2315,cstatus_csv_dumper_2315);
    fifo_csv_dumper_2316 = new("./depth2316.csv");
    cstatus_csv_dumper_2316 = new("./chan_status2316.csv");
    fifo_monitor_2316 = new(fifo_csv_dumper_2316,fifo_intf_2316,cstatus_csv_dumper_2316);
    fifo_csv_dumper_2317 = new("./depth2317.csv");
    cstatus_csv_dumper_2317 = new("./chan_status2317.csv");
    fifo_monitor_2317 = new(fifo_csv_dumper_2317,fifo_intf_2317,cstatus_csv_dumper_2317);
    fifo_csv_dumper_2318 = new("./depth2318.csv");
    cstatus_csv_dumper_2318 = new("./chan_status2318.csv");
    fifo_monitor_2318 = new(fifo_csv_dumper_2318,fifo_intf_2318,cstatus_csv_dumper_2318);
    fifo_csv_dumper_2319 = new("./depth2319.csv");
    cstatus_csv_dumper_2319 = new("./chan_status2319.csv");
    fifo_monitor_2319 = new(fifo_csv_dumper_2319,fifo_intf_2319,cstatus_csv_dumper_2319);
    fifo_csv_dumper_2320 = new("./depth2320.csv");
    cstatus_csv_dumper_2320 = new("./chan_status2320.csv");
    fifo_monitor_2320 = new(fifo_csv_dumper_2320,fifo_intf_2320,cstatus_csv_dumper_2320);
    fifo_csv_dumper_2321 = new("./depth2321.csv");
    cstatus_csv_dumper_2321 = new("./chan_status2321.csv");
    fifo_monitor_2321 = new(fifo_csv_dumper_2321,fifo_intf_2321,cstatus_csv_dumper_2321);
    fifo_csv_dumper_2322 = new("./depth2322.csv");
    cstatus_csv_dumper_2322 = new("./chan_status2322.csv");
    fifo_monitor_2322 = new(fifo_csv_dumper_2322,fifo_intf_2322,cstatus_csv_dumper_2322);
    fifo_csv_dumper_2323 = new("./depth2323.csv");
    cstatus_csv_dumper_2323 = new("./chan_status2323.csv");
    fifo_monitor_2323 = new(fifo_csv_dumper_2323,fifo_intf_2323,cstatus_csv_dumper_2323);
    fifo_csv_dumper_2324 = new("./depth2324.csv");
    cstatus_csv_dumper_2324 = new("./chan_status2324.csv");
    fifo_monitor_2324 = new(fifo_csv_dumper_2324,fifo_intf_2324,cstatus_csv_dumper_2324);
    fifo_csv_dumper_2325 = new("./depth2325.csv");
    cstatus_csv_dumper_2325 = new("./chan_status2325.csv");
    fifo_monitor_2325 = new(fifo_csv_dumper_2325,fifo_intf_2325,cstatus_csv_dumper_2325);
    fifo_csv_dumper_2326 = new("./depth2326.csv");
    cstatus_csv_dumper_2326 = new("./chan_status2326.csv");
    fifo_monitor_2326 = new(fifo_csv_dumper_2326,fifo_intf_2326,cstatus_csv_dumper_2326);
    fifo_csv_dumper_2327 = new("./depth2327.csv");
    cstatus_csv_dumper_2327 = new("./chan_status2327.csv");
    fifo_monitor_2327 = new(fifo_csv_dumper_2327,fifo_intf_2327,cstatus_csv_dumper_2327);
    fifo_csv_dumper_2328 = new("./depth2328.csv");
    cstatus_csv_dumper_2328 = new("./chan_status2328.csv");
    fifo_monitor_2328 = new(fifo_csv_dumper_2328,fifo_intf_2328,cstatus_csv_dumper_2328);
    fifo_csv_dumper_2329 = new("./depth2329.csv");
    cstatus_csv_dumper_2329 = new("./chan_status2329.csv");
    fifo_monitor_2329 = new(fifo_csv_dumper_2329,fifo_intf_2329,cstatus_csv_dumper_2329);
    fifo_csv_dumper_2330 = new("./depth2330.csv");
    cstatus_csv_dumper_2330 = new("./chan_status2330.csv");
    fifo_monitor_2330 = new(fifo_csv_dumper_2330,fifo_intf_2330,cstatus_csv_dumper_2330);
    fifo_csv_dumper_2331 = new("./depth2331.csv");
    cstatus_csv_dumper_2331 = new("./chan_status2331.csv");
    fifo_monitor_2331 = new(fifo_csv_dumper_2331,fifo_intf_2331,cstatus_csv_dumper_2331);
    fifo_csv_dumper_2332 = new("./depth2332.csv");
    cstatus_csv_dumper_2332 = new("./chan_status2332.csv");
    fifo_monitor_2332 = new(fifo_csv_dumper_2332,fifo_intf_2332,cstatus_csv_dumper_2332);
    fifo_csv_dumper_2333 = new("./depth2333.csv");
    cstatus_csv_dumper_2333 = new("./chan_status2333.csv");
    fifo_monitor_2333 = new(fifo_csv_dumper_2333,fifo_intf_2333,cstatus_csv_dumper_2333);
    fifo_csv_dumper_2334 = new("./depth2334.csv");
    cstatus_csv_dumper_2334 = new("./chan_status2334.csv");
    fifo_monitor_2334 = new(fifo_csv_dumper_2334,fifo_intf_2334,cstatus_csv_dumper_2334);
    fifo_csv_dumper_2335 = new("./depth2335.csv");
    cstatus_csv_dumper_2335 = new("./chan_status2335.csv");
    fifo_monitor_2335 = new(fifo_csv_dumper_2335,fifo_intf_2335,cstatus_csv_dumper_2335);
    fifo_csv_dumper_2336 = new("./depth2336.csv");
    cstatus_csv_dumper_2336 = new("./chan_status2336.csv");
    fifo_monitor_2336 = new(fifo_csv_dumper_2336,fifo_intf_2336,cstatus_csv_dumper_2336);
    fifo_csv_dumper_2337 = new("./depth2337.csv");
    cstatus_csv_dumper_2337 = new("./chan_status2337.csv");
    fifo_monitor_2337 = new(fifo_csv_dumper_2337,fifo_intf_2337,cstatus_csv_dumper_2337);
    fifo_csv_dumper_2338 = new("./depth2338.csv");
    cstatus_csv_dumper_2338 = new("./chan_status2338.csv");
    fifo_monitor_2338 = new(fifo_csv_dumper_2338,fifo_intf_2338,cstatus_csv_dumper_2338);
    fifo_csv_dumper_2339 = new("./depth2339.csv");
    cstatus_csv_dumper_2339 = new("./chan_status2339.csv");
    fifo_monitor_2339 = new(fifo_csv_dumper_2339,fifo_intf_2339,cstatus_csv_dumper_2339);
    fifo_csv_dumper_2340 = new("./depth2340.csv");
    cstatus_csv_dumper_2340 = new("./chan_status2340.csv");
    fifo_monitor_2340 = new(fifo_csv_dumper_2340,fifo_intf_2340,cstatus_csv_dumper_2340);
    fifo_csv_dumper_2341 = new("./depth2341.csv");
    cstatus_csv_dumper_2341 = new("./chan_status2341.csv");
    fifo_monitor_2341 = new(fifo_csv_dumper_2341,fifo_intf_2341,cstatus_csv_dumper_2341);
    fifo_csv_dumper_2342 = new("./depth2342.csv");
    cstatus_csv_dumper_2342 = new("./chan_status2342.csv");
    fifo_monitor_2342 = new(fifo_csv_dumper_2342,fifo_intf_2342,cstatus_csv_dumper_2342);
    fifo_csv_dumper_2343 = new("./depth2343.csv");
    cstatus_csv_dumper_2343 = new("./chan_status2343.csv");
    fifo_monitor_2343 = new(fifo_csv_dumper_2343,fifo_intf_2343,cstatus_csv_dumper_2343);
    fifo_csv_dumper_2344 = new("./depth2344.csv");
    cstatus_csv_dumper_2344 = new("./chan_status2344.csv");
    fifo_monitor_2344 = new(fifo_csv_dumper_2344,fifo_intf_2344,cstatus_csv_dumper_2344);
    fifo_csv_dumper_2345 = new("./depth2345.csv");
    cstatus_csv_dumper_2345 = new("./chan_status2345.csv");
    fifo_monitor_2345 = new(fifo_csv_dumper_2345,fifo_intf_2345,cstatus_csv_dumper_2345);
    fifo_csv_dumper_2346 = new("./depth2346.csv");
    cstatus_csv_dumper_2346 = new("./chan_status2346.csv");
    fifo_monitor_2346 = new(fifo_csv_dumper_2346,fifo_intf_2346,cstatus_csv_dumper_2346);
    fifo_csv_dumper_2347 = new("./depth2347.csv");
    cstatus_csv_dumper_2347 = new("./chan_status2347.csv");
    fifo_monitor_2347 = new(fifo_csv_dumper_2347,fifo_intf_2347,cstatus_csv_dumper_2347);
    fifo_csv_dumper_2348 = new("./depth2348.csv");
    cstatus_csv_dumper_2348 = new("./chan_status2348.csv");
    fifo_monitor_2348 = new(fifo_csv_dumper_2348,fifo_intf_2348,cstatus_csv_dumper_2348);
    fifo_csv_dumper_2349 = new("./depth2349.csv");
    cstatus_csv_dumper_2349 = new("./chan_status2349.csv");
    fifo_monitor_2349 = new(fifo_csv_dumper_2349,fifo_intf_2349,cstatus_csv_dumper_2349);
    fifo_csv_dumper_2350 = new("./depth2350.csv");
    cstatus_csv_dumper_2350 = new("./chan_status2350.csv");
    fifo_monitor_2350 = new(fifo_csv_dumper_2350,fifo_intf_2350,cstatus_csv_dumper_2350);
    fifo_csv_dumper_2351 = new("./depth2351.csv");
    cstatus_csv_dumper_2351 = new("./chan_status2351.csv");
    fifo_monitor_2351 = new(fifo_csv_dumper_2351,fifo_intf_2351,cstatus_csv_dumper_2351);
    fifo_csv_dumper_2352 = new("./depth2352.csv");
    cstatus_csv_dumper_2352 = new("./chan_status2352.csv");
    fifo_monitor_2352 = new(fifo_csv_dumper_2352,fifo_intf_2352,cstatus_csv_dumper_2352);
    fifo_csv_dumper_2353 = new("./depth2353.csv");
    cstatus_csv_dumper_2353 = new("./chan_status2353.csv");
    fifo_monitor_2353 = new(fifo_csv_dumper_2353,fifo_intf_2353,cstatus_csv_dumper_2353);
    fifo_csv_dumper_2354 = new("./depth2354.csv");
    cstatus_csv_dumper_2354 = new("./chan_status2354.csv");
    fifo_monitor_2354 = new(fifo_csv_dumper_2354,fifo_intf_2354,cstatus_csv_dumper_2354);
    fifo_csv_dumper_2355 = new("./depth2355.csv");
    cstatus_csv_dumper_2355 = new("./chan_status2355.csv");
    fifo_monitor_2355 = new(fifo_csv_dumper_2355,fifo_intf_2355,cstatus_csv_dumper_2355);
    fifo_csv_dumper_2356 = new("./depth2356.csv");
    cstatus_csv_dumper_2356 = new("./chan_status2356.csv");
    fifo_monitor_2356 = new(fifo_csv_dumper_2356,fifo_intf_2356,cstatus_csv_dumper_2356);
    fifo_csv_dumper_2357 = new("./depth2357.csv");
    cstatus_csv_dumper_2357 = new("./chan_status2357.csv");
    fifo_monitor_2357 = new(fifo_csv_dumper_2357,fifo_intf_2357,cstatus_csv_dumper_2357);
    fifo_csv_dumper_2358 = new("./depth2358.csv");
    cstatus_csv_dumper_2358 = new("./chan_status2358.csv");
    fifo_monitor_2358 = new(fifo_csv_dumper_2358,fifo_intf_2358,cstatus_csv_dumper_2358);
    fifo_csv_dumper_2359 = new("./depth2359.csv");
    cstatus_csv_dumper_2359 = new("./chan_status2359.csv");
    fifo_monitor_2359 = new(fifo_csv_dumper_2359,fifo_intf_2359,cstatus_csv_dumper_2359);
    fifo_csv_dumper_2360 = new("./depth2360.csv");
    cstatus_csv_dumper_2360 = new("./chan_status2360.csv");
    fifo_monitor_2360 = new(fifo_csv_dumper_2360,fifo_intf_2360,cstatus_csv_dumper_2360);
    fifo_csv_dumper_2361 = new("./depth2361.csv");
    cstatus_csv_dumper_2361 = new("./chan_status2361.csv");
    fifo_monitor_2361 = new(fifo_csv_dumper_2361,fifo_intf_2361,cstatus_csv_dumper_2361);
    fifo_csv_dumper_2362 = new("./depth2362.csv");
    cstatus_csv_dumper_2362 = new("./chan_status2362.csv");
    fifo_monitor_2362 = new(fifo_csv_dumper_2362,fifo_intf_2362,cstatus_csv_dumper_2362);
    fifo_csv_dumper_2363 = new("./depth2363.csv");
    cstatus_csv_dumper_2363 = new("./chan_status2363.csv");
    fifo_monitor_2363 = new(fifo_csv_dumper_2363,fifo_intf_2363,cstatus_csv_dumper_2363);
    fifo_csv_dumper_2364 = new("./depth2364.csv");
    cstatus_csv_dumper_2364 = new("./chan_status2364.csv");
    fifo_monitor_2364 = new(fifo_csv_dumper_2364,fifo_intf_2364,cstatus_csv_dumper_2364);
    fifo_csv_dumper_2365 = new("./depth2365.csv");
    cstatus_csv_dumper_2365 = new("./chan_status2365.csv");
    fifo_monitor_2365 = new(fifo_csv_dumper_2365,fifo_intf_2365,cstatus_csv_dumper_2365);
    fifo_csv_dumper_2366 = new("./depth2366.csv");
    cstatus_csv_dumper_2366 = new("./chan_status2366.csv");
    fifo_monitor_2366 = new(fifo_csv_dumper_2366,fifo_intf_2366,cstatus_csv_dumper_2366);
    fifo_csv_dumper_2367 = new("./depth2367.csv");
    cstatus_csv_dumper_2367 = new("./chan_status2367.csv");
    fifo_monitor_2367 = new(fifo_csv_dumper_2367,fifo_intf_2367,cstatus_csv_dumper_2367);
    fifo_csv_dumper_2368 = new("./depth2368.csv");
    cstatus_csv_dumper_2368 = new("./chan_status2368.csv");
    fifo_monitor_2368 = new(fifo_csv_dumper_2368,fifo_intf_2368,cstatus_csv_dumper_2368);
    fifo_csv_dumper_2369 = new("./depth2369.csv");
    cstatus_csv_dumper_2369 = new("./chan_status2369.csv");
    fifo_monitor_2369 = new(fifo_csv_dumper_2369,fifo_intf_2369,cstatus_csv_dumper_2369);
    fifo_csv_dumper_2370 = new("./depth2370.csv");
    cstatus_csv_dumper_2370 = new("./chan_status2370.csv");
    fifo_monitor_2370 = new(fifo_csv_dumper_2370,fifo_intf_2370,cstatus_csv_dumper_2370);
    fifo_csv_dumper_2371 = new("./depth2371.csv");
    cstatus_csv_dumper_2371 = new("./chan_status2371.csv");
    fifo_monitor_2371 = new(fifo_csv_dumper_2371,fifo_intf_2371,cstatus_csv_dumper_2371);
    fifo_csv_dumper_2372 = new("./depth2372.csv");
    cstatus_csv_dumper_2372 = new("./chan_status2372.csv");
    fifo_monitor_2372 = new(fifo_csv_dumper_2372,fifo_intf_2372,cstatus_csv_dumper_2372);
    fifo_csv_dumper_2373 = new("./depth2373.csv");
    cstatus_csv_dumper_2373 = new("./chan_status2373.csv");
    fifo_monitor_2373 = new(fifo_csv_dumper_2373,fifo_intf_2373,cstatus_csv_dumper_2373);
    fifo_csv_dumper_2374 = new("./depth2374.csv");
    cstatus_csv_dumper_2374 = new("./chan_status2374.csv");
    fifo_monitor_2374 = new(fifo_csv_dumper_2374,fifo_intf_2374,cstatus_csv_dumper_2374);
    fifo_csv_dumper_2375 = new("./depth2375.csv");
    cstatus_csv_dumper_2375 = new("./chan_status2375.csv");
    fifo_monitor_2375 = new(fifo_csv_dumper_2375,fifo_intf_2375,cstatus_csv_dumper_2375);
    fifo_csv_dumper_2376 = new("./depth2376.csv");
    cstatus_csv_dumper_2376 = new("./chan_status2376.csv");
    fifo_monitor_2376 = new(fifo_csv_dumper_2376,fifo_intf_2376,cstatus_csv_dumper_2376);
    fifo_csv_dumper_2377 = new("./depth2377.csv");
    cstatus_csv_dumper_2377 = new("./chan_status2377.csv");
    fifo_monitor_2377 = new(fifo_csv_dumper_2377,fifo_intf_2377,cstatus_csv_dumper_2377);
    fifo_csv_dumper_2378 = new("./depth2378.csv");
    cstatus_csv_dumper_2378 = new("./chan_status2378.csv");
    fifo_monitor_2378 = new(fifo_csv_dumper_2378,fifo_intf_2378,cstatus_csv_dumper_2378);
    fifo_csv_dumper_2379 = new("./depth2379.csv");
    cstatus_csv_dumper_2379 = new("./chan_status2379.csv");
    fifo_monitor_2379 = new(fifo_csv_dumper_2379,fifo_intf_2379,cstatus_csv_dumper_2379);
    fifo_csv_dumper_2380 = new("./depth2380.csv");
    cstatus_csv_dumper_2380 = new("./chan_status2380.csv");
    fifo_monitor_2380 = new(fifo_csv_dumper_2380,fifo_intf_2380,cstatus_csv_dumper_2380);
    fifo_csv_dumper_2381 = new("./depth2381.csv");
    cstatus_csv_dumper_2381 = new("./chan_status2381.csv");
    fifo_monitor_2381 = new(fifo_csv_dumper_2381,fifo_intf_2381,cstatus_csv_dumper_2381);
    fifo_csv_dumper_2382 = new("./depth2382.csv");
    cstatus_csv_dumper_2382 = new("./chan_status2382.csv");
    fifo_monitor_2382 = new(fifo_csv_dumper_2382,fifo_intf_2382,cstatus_csv_dumper_2382);
    fifo_csv_dumper_2383 = new("./depth2383.csv");
    cstatus_csv_dumper_2383 = new("./chan_status2383.csv");
    fifo_monitor_2383 = new(fifo_csv_dumper_2383,fifo_intf_2383,cstatus_csv_dumper_2383);
    fifo_csv_dumper_2384 = new("./depth2384.csv");
    cstatus_csv_dumper_2384 = new("./chan_status2384.csv");
    fifo_monitor_2384 = new(fifo_csv_dumper_2384,fifo_intf_2384,cstatus_csv_dumper_2384);
    fifo_csv_dumper_2385 = new("./depth2385.csv");
    cstatus_csv_dumper_2385 = new("./chan_status2385.csv");
    fifo_monitor_2385 = new(fifo_csv_dumper_2385,fifo_intf_2385,cstatus_csv_dumper_2385);
    fifo_csv_dumper_2386 = new("./depth2386.csv");
    cstatus_csv_dumper_2386 = new("./chan_status2386.csv");
    fifo_monitor_2386 = new(fifo_csv_dumper_2386,fifo_intf_2386,cstatus_csv_dumper_2386);
    fifo_csv_dumper_2387 = new("./depth2387.csv");
    cstatus_csv_dumper_2387 = new("./chan_status2387.csv");
    fifo_monitor_2387 = new(fifo_csv_dumper_2387,fifo_intf_2387,cstatus_csv_dumper_2387);
    fifo_csv_dumper_2388 = new("./depth2388.csv");
    cstatus_csv_dumper_2388 = new("./chan_status2388.csv");
    fifo_monitor_2388 = new(fifo_csv_dumper_2388,fifo_intf_2388,cstatus_csv_dumper_2388);
    fifo_csv_dumper_2389 = new("./depth2389.csv");
    cstatus_csv_dumper_2389 = new("./chan_status2389.csv");
    fifo_monitor_2389 = new(fifo_csv_dumper_2389,fifo_intf_2389,cstatus_csv_dumper_2389);
    fifo_csv_dumper_2390 = new("./depth2390.csv");
    cstatus_csv_dumper_2390 = new("./chan_status2390.csv");
    fifo_monitor_2390 = new(fifo_csv_dumper_2390,fifo_intf_2390,cstatus_csv_dumper_2390);
    fifo_csv_dumper_2391 = new("./depth2391.csv");
    cstatus_csv_dumper_2391 = new("./chan_status2391.csv");
    fifo_monitor_2391 = new(fifo_csv_dumper_2391,fifo_intf_2391,cstatus_csv_dumper_2391);
    fifo_csv_dumper_2392 = new("./depth2392.csv");
    cstatus_csv_dumper_2392 = new("./chan_status2392.csv");
    fifo_monitor_2392 = new(fifo_csv_dumper_2392,fifo_intf_2392,cstatus_csv_dumper_2392);
    fifo_csv_dumper_2393 = new("./depth2393.csv");
    cstatus_csv_dumper_2393 = new("./chan_status2393.csv");
    fifo_monitor_2393 = new(fifo_csv_dumper_2393,fifo_intf_2393,cstatus_csv_dumper_2393);
    fifo_csv_dumper_2394 = new("./depth2394.csv");
    cstatus_csv_dumper_2394 = new("./chan_status2394.csv");
    fifo_monitor_2394 = new(fifo_csv_dumper_2394,fifo_intf_2394,cstatus_csv_dumper_2394);
    fifo_csv_dumper_2395 = new("./depth2395.csv");
    cstatus_csv_dumper_2395 = new("./chan_status2395.csv");
    fifo_monitor_2395 = new(fifo_csv_dumper_2395,fifo_intf_2395,cstatus_csv_dumper_2395);
    fifo_csv_dumper_2396 = new("./depth2396.csv");
    cstatus_csv_dumper_2396 = new("./chan_status2396.csv");
    fifo_monitor_2396 = new(fifo_csv_dumper_2396,fifo_intf_2396,cstatus_csv_dumper_2396);
    fifo_csv_dumper_2397 = new("./depth2397.csv");
    cstatus_csv_dumper_2397 = new("./chan_status2397.csv");
    fifo_monitor_2397 = new(fifo_csv_dumper_2397,fifo_intf_2397,cstatus_csv_dumper_2397);
    fifo_csv_dumper_2398 = new("./depth2398.csv");
    cstatus_csv_dumper_2398 = new("./chan_status2398.csv");
    fifo_monitor_2398 = new(fifo_csv_dumper_2398,fifo_intf_2398,cstatus_csv_dumper_2398);
    fifo_csv_dumper_2399 = new("./depth2399.csv");
    cstatus_csv_dumper_2399 = new("./chan_status2399.csv");
    fifo_monitor_2399 = new(fifo_csv_dumper_2399,fifo_intf_2399,cstatus_csv_dumper_2399);
    fifo_csv_dumper_2400 = new("./depth2400.csv");
    cstatus_csv_dumper_2400 = new("./chan_status2400.csv");
    fifo_monitor_2400 = new(fifo_csv_dumper_2400,fifo_intf_2400,cstatus_csv_dumper_2400);
    fifo_csv_dumper_2401 = new("./depth2401.csv");
    cstatus_csv_dumper_2401 = new("./chan_status2401.csv");
    fifo_monitor_2401 = new(fifo_csv_dumper_2401,fifo_intf_2401,cstatus_csv_dumper_2401);
    fifo_csv_dumper_2402 = new("./depth2402.csv");
    cstatus_csv_dumper_2402 = new("./chan_status2402.csv");
    fifo_monitor_2402 = new(fifo_csv_dumper_2402,fifo_intf_2402,cstatus_csv_dumper_2402);
    fifo_csv_dumper_2403 = new("./depth2403.csv");
    cstatus_csv_dumper_2403 = new("./chan_status2403.csv");
    fifo_monitor_2403 = new(fifo_csv_dumper_2403,fifo_intf_2403,cstatus_csv_dumper_2403);
    fifo_csv_dumper_2404 = new("./depth2404.csv");
    cstatus_csv_dumper_2404 = new("./chan_status2404.csv");
    fifo_monitor_2404 = new(fifo_csv_dumper_2404,fifo_intf_2404,cstatus_csv_dumper_2404);
    fifo_csv_dumper_2405 = new("./depth2405.csv");
    cstatus_csv_dumper_2405 = new("./chan_status2405.csv");
    fifo_monitor_2405 = new(fifo_csv_dumper_2405,fifo_intf_2405,cstatus_csv_dumper_2405);
    fifo_csv_dumper_2406 = new("./depth2406.csv");
    cstatus_csv_dumper_2406 = new("./chan_status2406.csv");
    fifo_monitor_2406 = new(fifo_csv_dumper_2406,fifo_intf_2406,cstatus_csv_dumper_2406);
    fifo_csv_dumper_2407 = new("./depth2407.csv");
    cstatus_csv_dumper_2407 = new("./chan_status2407.csv");
    fifo_monitor_2407 = new(fifo_csv_dumper_2407,fifo_intf_2407,cstatus_csv_dumper_2407);
    fifo_csv_dumper_2408 = new("./depth2408.csv");
    cstatus_csv_dumper_2408 = new("./chan_status2408.csv");
    fifo_monitor_2408 = new(fifo_csv_dumper_2408,fifo_intf_2408,cstatus_csv_dumper_2408);
    fifo_csv_dumper_2409 = new("./depth2409.csv");
    cstatus_csv_dumper_2409 = new("./chan_status2409.csv");
    fifo_monitor_2409 = new(fifo_csv_dumper_2409,fifo_intf_2409,cstatus_csv_dumper_2409);
    fifo_csv_dumper_2410 = new("./depth2410.csv");
    cstatus_csv_dumper_2410 = new("./chan_status2410.csv");
    fifo_monitor_2410 = new(fifo_csv_dumper_2410,fifo_intf_2410,cstatus_csv_dumper_2410);
    fifo_csv_dumper_2411 = new("./depth2411.csv");
    cstatus_csv_dumper_2411 = new("./chan_status2411.csv");
    fifo_monitor_2411 = new(fifo_csv_dumper_2411,fifo_intf_2411,cstatus_csv_dumper_2411);
    fifo_csv_dumper_2412 = new("./depth2412.csv");
    cstatus_csv_dumper_2412 = new("./chan_status2412.csv");
    fifo_monitor_2412 = new(fifo_csv_dumper_2412,fifo_intf_2412,cstatus_csv_dumper_2412);
    fifo_csv_dumper_2413 = new("./depth2413.csv");
    cstatus_csv_dumper_2413 = new("./chan_status2413.csv");
    fifo_monitor_2413 = new(fifo_csv_dumper_2413,fifo_intf_2413,cstatus_csv_dumper_2413);
    fifo_csv_dumper_2414 = new("./depth2414.csv");
    cstatus_csv_dumper_2414 = new("./chan_status2414.csv");
    fifo_monitor_2414 = new(fifo_csv_dumper_2414,fifo_intf_2414,cstatus_csv_dumper_2414);
    fifo_csv_dumper_2415 = new("./depth2415.csv");
    cstatus_csv_dumper_2415 = new("./chan_status2415.csv");
    fifo_monitor_2415 = new(fifo_csv_dumper_2415,fifo_intf_2415,cstatus_csv_dumper_2415);
    fifo_csv_dumper_2416 = new("./depth2416.csv");
    cstatus_csv_dumper_2416 = new("./chan_status2416.csv");
    fifo_monitor_2416 = new(fifo_csv_dumper_2416,fifo_intf_2416,cstatus_csv_dumper_2416);
    fifo_csv_dumper_2417 = new("./depth2417.csv");
    cstatus_csv_dumper_2417 = new("./chan_status2417.csv");
    fifo_monitor_2417 = new(fifo_csv_dumper_2417,fifo_intf_2417,cstatus_csv_dumper_2417);
    fifo_csv_dumper_2418 = new("./depth2418.csv");
    cstatus_csv_dumper_2418 = new("./chan_status2418.csv");
    fifo_monitor_2418 = new(fifo_csv_dumper_2418,fifo_intf_2418,cstatus_csv_dumper_2418);
    fifo_csv_dumper_2419 = new("./depth2419.csv");
    cstatus_csv_dumper_2419 = new("./chan_status2419.csv");
    fifo_monitor_2419 = new(fifo_csv_dumper_2419,fifo_intf_2419,cstatus_csv_dumper_2419);
    fifo_csv_dumper_2420 = new("./depth2420.csv");
    cstatus_csv_dumper_2420 = new("./chan_status2420.csv");
    fifo_monitor_2420 = new(fifo_csv_dumper_2420,fifo_intf_2420,cstatus_csv_dumper_2420);
    fifo_csv_dumper_2421 = new("./depth2421.csv");
    cstatus_csv_dumper_2421 = new("./chan_status2421.csv");
    fifo_monitor_2421 = new(fifo_csv_dumper_2421,fifo_intf_2421,cstatus_csv_dumper_2421);
    fifo_csv_dumper_2422 = new("./depth2422.csv");
    cstatus_csv_dumper_2422 = new("./chan_status2422.csv");
    fifo_monitor_2422 = new(fifo_csv_dumper_2422,fifo_intf_2422,cstatus_csv_dumper_2422);
    fifo_csv_dumper_2423 = new("./depth2423.csv");
    cstatus_csv_dumper_2423 = new("./chan_status2423.csv");
    fifo_monitor_2423 = new(fifo_csv_dumper_2423,fifo_intf_2423,cstatus_csv_dumper_2423);
    fifo_csv_dumper_2424 = new("./depth2424.csv");
    cstatus_csv_dumper_2424 = new("./chan_status2424.csv");
    fifo_monitor_2424 = new(fifo_csv_dumper_2424,fifo_intf_2424,cstatus_csv_dumper_2424);
    fifo_csv_dumper_2425 = new("./depth2425.csv");
    cstatus_csv_dumper_2425 = new("./chan_status2425.csv");
    fifo_monitor_2425 = new(fifo_csv_dumper_2425,fifo_intf_2425,cstatus_csv_dumper_2425);
    fifo_csv_dumper_2426 = new("./depth2426.csv");
    cstatus_csv_dumper_2426 = new("./chan_status2426.csv");
    fifo_monitor_2426 = new(fifo_csv_dumper_2426,fifo_intf_2426,cstatus_csv_dumper_2426);
    fifo_csv_dumper_2427 = new("./depth2427.csv");
    cstatus_csv_dumper_2427 = new("./chan_status2427.csv");
    fifo_monitor_2427 = new(fifo_csv_dumper_2427,fifo_intf_2427,cstatus_csv_dumper_2427);
    fifo_csv_dumper_2428 = new("./depth2428.csv");
    cstatus_csv_dumper_2428 = new("./chan_status2428.csv");
    fifo_monitor_2428 = new(fifo_csv_dumper_2428,fifo_intf_2428,cstatus_csv_dumper_2428);
    fifo_csv_dumper_2429 = new("./depth2429.csv");
    cstatus_csv_dumper_2429 = new("./chan_status2429.csv");
    fifo_monitor_2429 = new(fifo_csv_dumper_2429,fifo_intf_2429,cstatus_csv_dumper_2429);
    fifo_csv_dumper_2430 = new("./depth2430.csv");
    cstatus_csv_dumper_2430 = new("./chan_status2430.csv");
    fifo_monitor_2430 = new(fifo_csv_dumper_2430,fifo_intf_2430,cstatus_csv_dumper_2430);
    fifo_csv_dumper_2431 = new("./depth2431.csv");
    cstatus_csv_dumper_2431 = new("./chan_status2431.csv");
    fifo_monitor_2431 = new(fifo_csv_dumper_2431,fifo_intf_2431,cstatus_csv_dumper_2431);
    fifo_csv_dumper_2432 = new("./depth2432.csv");
    cstatus_csv_dumper_2432 = new("./chan_status2432.csv");
    fifo_monitor_2432 = new(fifo_csv_dumper_2432,fifo_intf_2432,cstatus_csv_dumper_2432);
    fifo_csv_dumper_2433 = new("./depth2433.csv");
    cstatus_csv_dumper_2433 = new("./chan_status2433.csv");
    fifo_monitor_2433 = new(fifo_csv_dumper_2433,fifo_intf_2433,cstatus_csv_dumper_2433);
    fifo_csv_dumper_2434 = new("./depth2434.csv");
    cstatus_csv_dumper_2434 = new("./chan_status2434.csv");
    fifo_monitor_2434 = new(fifo_csv_dumper_2434,fifo_intf_2434,cstatus_csv_dumper_2434);
    fifo_csv_dumper_2435 = new("./depth2435.csv");
    cstatus_csv_dumper_2435 = new("./chan_status2435.csv");
    fifo_monitor_2435 = new(fifo_csv_dumper_2435,fifo_intf_2435,cstatus_csv_dumper_2435);
    fifo_csv_dumper_2436 = new("./depth2436.csv");
    cstatus_csv_dumper_2436 = new("./chan_status2436.csv");
    fifo_monitor_2436 = new(fifo_csv_dumper_2436,fifo_intf_2436,cstatus_csv_dumper_2436);
    fifo_csv_dumper_2437 = new("./depth2437.csv");
    cstatus_csv_dumper_2437 = new("./chan_status2437.csv");
    fifo_monitor_2437 = new(fifo_csv_dumper_2437,fifo_intf_2437,cstatus_csv_dumper_2437);
    fifo_csv_dumper_2438 = new("./depth2438.csv");
    cstatus_csv_dumper_2438 = new("./chan_status2438.csv");
    fifo_monitor_2438 = new(fifo_csv_dumper_2438,fifo_intf_2438,cstatus_csv_dumper_2438);
    fifo_csv_dumper_2439 = new("./depth2439.csv");
    cstatus_csv_dumper_2439 = new("./chan_status2439.csv");
    fifo_monitor_2439 = new(fifo_csv_dumper_2439,fifo_intf_2439,cstatus_csv_dumper_2439);
    fifo_csv_dumper_2440 = new("./depth2440.csv");
    cstatus_csv_dumper_2440 = new("./chan_status2440.csv");
    fifo_monitor_2440 = new(fifo_csv_dumper_2440,fifo_intf_2440,cstatus_csv_dumper_2440);
    fifo_csv_dumper_2441 = new("./depth2441.csv");
    cstatus_csv_dumper_2441 = new("./chan_status2441.csv");
    fifo_monitor_2441 = new(fifo_csv_dumper_2441,fifo_intf_2441,cstatus_csv_dumper_2441);
    fifo_csv_dumper_2442 = new("./depth2442.csv");
    cstatus_csv_dumper_2442 = new("./chan_status2442.csv");
    fifo_monitor_2442 = new(fifo_csv_dumper_2442,fifo_intf_2442,cstatus_csv_dumper_2442);
    fifo_csv_dumper_2443 = new("./depth2443.csv");
    cstatus_csv_dumper_2443 = new("./chan_status2443.csv");
    fifo_monitor_2443 = new(fifo_csv_dumper_2443,fifo_intf_2443,cstatus_csv_dumper_2443);
    fifo_csv_dumper_2444 = new("./depth2444.csv");
    cstatus_csv_dumper_2444 = new("./chan_status2444.csv");
    fifo_monitor_2444 = new(fifo_csv_dumper_2444,fifo_intf_2444,cstatus_csv_dumper_2444);
    fifo_csv_dumper_2445 = new("./depth2445.csv");
    cstatus_csv_dumper_2445 = new("./chan_status2445.csv");
    fifo_monitor_2445 = new(fifo_csv_dumper_2445,fifo_intf_2445,cstatus_csv_dumper_2445);
    fifo_csv_dumper_2446 = new("./depth2446.csv");
    cstatus_csv_dumper_2446 = new("./chan_status2446.csv");
    fifo_monitor_2446 = new(fifo_csv_dumper_2446,fifo_intf_2446,cstatus_csv_dumper_2446);
    fifo_csv_dumper_2447 = new("./depth2447.csv");
    cstatus_csv_dumper_2447 = new("./chan_status2447.csv");
    fifo_monitor_2447 = new(fifo_csv_dumper_2447,fifo_intf_2447,cstatus_csv_dumper_2447);
    fifo_csv_dumper_2448 = new("./depth2448.csv");
    cstatus_csv_dumper_2448 = new("./chan_status2448.csv");
    fifo_monitor_2448 = new(fifo_csv_dumper_2448,fifo_intf_2448,cstatus_csv_dumper_2448);
    fifo_csv_dumper_2449 = new("./depth2449.csv");
    cstatus_csv_dumper_2449 = new("./chan_status2449.csv");
    fifo_monitor_2449 = new(fifo_csv_dumper_2449,fifo_intf_2449,cstatus_csv_dumper_2449);
    fifo_csv_dumper_2450 = new("./depth2450.csv");
    cstatus_csv_dumper_2450 = new("./chan_status2450.csv");
    fifo_monitor_2450 = new(fifo_csv_dumper_2450,fifo_intf_2450,cstatus_csv_dumper_2450);
    fifo_csv_dumper_2451 = new("./depth2451.csv");
    cstatus_csv_dumper_2451 = new("./chan_status2451.csv");
    fifo_monitor_2451 = new(fifo_csv_dumper_2451,fifo_intf_2451,cstatus_csv_dumper_2451);
    fifo_csv_dumper_2452 = new("./depth2452.csv");
    cstatus_csv_dumper_2452 = new("./chan_status2452.csv");
    fifo_monitor_2452 = new(fifo_csv_dumper_2452,fifo_intf_2452,cstatus_csv_dumper_2452);
    fifo_csv_dumper_2453 = new("./depth2453.csv");
    cstatus_csv_dumper_2453 = new("./chan_status2453.csv");
    fifo_monitor_2453 = new(fifo_csv_dumper_2453,fifo_intf_2453,cstatus_csv_dumper_2453);
    fifo_csv_dumper_2454 = new("./depth2454.csv");
    cstatus_csv_dumper_2454 = new("./chan_status2454.csv");
    fifo_monitor_2454 = new(fifo_csv_dumper_2454,fifo_intf_2454,cstatus_csv_dumper_2454);
    fifo_csv_dumper_2455 = new("./depth2455.csv");
    cstatus_csv_dumper_2455 = new("./chan_status2455.csv");
    fifo_monitor_2455 = new(fifo_csv_dumper_2455,fifo_intf_2455,cstatus_csv_dumper_2455);
    fifo_csv_dumper_2456 = new("./depth2456.csv");
    cstatus_csv_dumper_2456 = new("./chan_status2456.csv");
    fifo_monitor_2456 = new(fifo_csv_dumper_2456,fifo_intf_2456,cstatus_csv_dumper_2456);
    fifo_csv_dumper_2457 = new("./depth2457.csv");
    cstatus_csv_dumper_2457 = new("./chan_status2457.csv");
    fifo_monitor_2457 = new(fifo_csv_dumper_2457,fifo_intf_2457,cstatus_csv_dumper_2457);
    fifo_csv_dumper_2458 = new("./depth2458.csv");
    cstatus_csv_dumper_2458 = new("./chan_status2458.csv");
    fifo_monitor_2458 = new(fifo_csv_dumper_2458,fifo_intf_2458,cstatus_csv_dumper_2458);
    fifo_csv_dumper_2459 = new("./depth2459.csv");
    cstatus_csv_dumper_2459 = new("./chan_status2459.csv");
    fifo_monitor_2459 = new(fifo_csv_dumper_2459,fifo_intf_2459,cstatus_csv_dumper_2459);
    fifo_csv_dumper_2460 = new("./depth2460.csv");
    cstatus_csv_dumper_2460 = new("./chan_status2460.csv");
    fifo_monitor_2460 = new(fifo_csv_dumper_2460,fifo_intf_2460,cstatus_csv_dumper_2460);
    fifo_csv_dumper_2461 = new("./depth2461.csv");
    cstatus_csv_dumper_2461 = new("./chan_status2461.csv");
    fifo_monitor_2461 = new(fifo_csv_dumper_2461,fifo_intf_2461,cstatus_csv_dumper_2461);
    fifo_csv_dumper_2462 = new("./depth2462.csv");
    cstatus_csv_dumper_2462 = new("./chan_status2462.csv");
    fifo_monitor_2462 = new(fifo_csv_dumper_2462,fifo_intf_2462,cstatus_csv_dumper_2462);
    fifo_csv_dumper_2463 = new("./depth2463.csv");
    cstatus_csv_dumper_2463 = new("./chan_status2463.csv");
    fifo_monitor_2463 = new(fifo_csv_dumper_2463,fifo_intf_2463,cstatus_csv_dumper_2463);
    fifo_csv_dumper_2464 = new("./depth2464.csv");
    cstatus_csv_dumper_2464 = new("./chan_status2464.csv");
    fifo_monitor_2464 = new(fifo_csv_dumper_2464,fifo_intf_2464,cstatus_csv_dumper_2464);
    fifo_csv_dumper_2465 = new("./depth2465.csv");
    cstatus_csv_dumper_2465 = new("./chan_status2465.csv");
    fifo_monitor_2465 = new(fifo_csv_dumper_2465,fifo_intf_2465,cstatus_csv_dumper_2465);
    fifo_csv_dumper_2466 = new("./depth2466.csv");
    cstatus_csv_dumper_2466 = new("./chan_status2466.csv");
    fifo_monitor_2466 = new(fifo_csv_dumper_2466,fifo_intf_2466,cstatus_csv_dumper_2466);
    fifo_csv_dumper_2467 = new("./depth2467.csv");
    cstatus_csv_dumper_2467 = new("./chan_status2467.csv");
    fifo_monitor_2467 = new(fifo_csv_dumper_2467,fifo_intf_2467,cstatus_csv_dumper_2467);
    fifo_csv_dumper_2468 = new("./depth2468.csv");
    cstatus_csv_dumper_2468 = new("./chan_status2468.csv");
    fifo_monitor_2468 = new(fifo_csv_dumper_2468,fifo_intf_2468,cstatus_csv_dumper_2468);
    fifo_csv_dumper_2469 = new("./depth2469.csv");
    cstatus_csv_dumper_2469 = new("./chan_status2469.csv");
    fifo_monitor_2469 = new(fifo_csv_dumper_2469,fifo_intf_2469,cstatus_csv_dumper_2469);
    fifo_csv_dumper_2470 = new("./depth2470.csv");
    cstatus_csv_dumper_2470 = new("./chan_status2470.csv");
    fifo_monitor_2470 = new(fifo_csv_dumper_2470,fifo_intf_2470,cstatus_csv_dumper_2470);
    fifo_csv_dumper_2471 = new("./depth2471.csv");
    cstatus_csv_dumper_2471 = new("./chan_status2471.csv");
    fifo_monitor_2471 = new(fifo_csv_dumper_2471,fifo_intf_2471,cstatus_csv_dumper_2471);
    fifo_csv_dumper_2472 = new("./depth2472.csv");
    cstatus_csv_dumper_2472 = new("./chan_status2472.csv");
    fifo_monitor_2472 = new(fifo_csv_dumper_2472,fifo_intf_2472,cstatus_csv_dumper_2472);
    fifo_csv_dumper_2473 = new("./depth2473.csv");
    cstatus_csv_dumper_2473 = new("./chan_status2473.csv");
    fifo_monitor_2473 = new(fifo_csv_dumper_2473,fifo_intf_2473,cstatus_csv_dumper_2473);
    fifo_csv_dumper_2474 = new("./depth2474.csv");
    cstatus_csv_dumper_2474 = new("./chan_status2474.csv");
    fifo_monitor_2474 = new(fifo_csv_dumper_2474,fifo_intf_2474,cstatus_csv_dumper_2474);
    fifo_csv_dumper_2475 = new("./depth2475.csv");
    cstatus_csv_dumper_2475 = new("./chan_status2475.csv");
    fifo_monitor_2475 = new(fifo_csv_dumper_2475,fifo_intf_2475,cstatus_csv_dumper_2475);
    fifo_csv_dumper_2476 = new("./depth2476.csv");
    cstatus_csv_dumper_2476 = new("./chan_status2476.csv");
    fifo_monitor_2476 = new(fifo_csv_dumper_2476,fifo_intf_2476,cstatus_csv_dumper_2476);
    fifo_csv_dumper_2477 = new("./depth2477.csv");
    cstatus_csv_dumper_2477 = new("./chan_status2477.csv");
    fifo_monitor_2477 = new(fifo_csv_dumper_2477,fifo_intf_2477,cstatus_csv_dumper_2477);
    fifo_csv_dumper_2478 = new("./depth2478.csv");
    cstatus_csv_dumper_2478 = new("./chan_status2478.csv");
    fifo_monitor_2478 = new(fifo_csv_dumper_2478,fifo_intf_2478,cstatus_csv_dumper_2478);
    fifo_csv_dumper_2479 = new("./depth2479.csv");
    cstatus_csv_dumper_2479 = new("./chan_status2479.csv");
    fifo_monitor_2479 = new(fifo_csv_dumper_2479,fifo_intf_2479,cstatus_csv_dumper_2479);
    fifo_csv_dumper_2480 = new("./depth2480.csv");
    cstatus_csv_dumper_2480 = new("./chan_status2480.csv");
    fifo_monitor_2480 = new(fifo_csv_dumper_2480,fifo_intf_2480,cstatus_csv_dumper_2480);
    fifo_csv_dumper_2481 = new("./depth2481.csv");
    cstatus_csv_dumper_2481 = new("./chan_status2481.csv");
    fifo_monitor_2481 = new(fifo_csv_dumper_2481,fifo_intf_2481,cstatus_csv_dumper_2481);
    fifo_csv_dumper_2482 = new("./depth2482.csv");
    cstatus_csv_dumper_2482 = new("./chan_status2482.csv");
    fifo_monitor_2482 = new(fifo_csv_dumper_2482,fifo_intf_2482,cstatus_csv_dumper_2482);
    fifo_csv_dumper_2483 = new("./depth2483.csv");
    cstatus_csv_dumper_2483 = new("./chan_status2483.csv");
    fifo_monitor_2483 = new(fifo_csv_dumper_2483,fifo_intf_2483,cstatus_csv_dumper_2483);
    fifo_csv_dumper_2484 = new("./depth2484.csv");
    cstatus_csv_dumper_2484 = new("./chan_status2484.csv");
    fifo_monitor_2484 = new(fifo_csv_dumper_2484,fifo_intf_2484,cstatus_csv_dumper_2484);
    fifo_csv_dumper_2485 = new("./depth2485.csv");
    cstatus_csv_dumper_2485 = new("./chan_status2485.csv");
    fifo_monitor_2485 = new(fifo_csv_dumper_2485,fifo_intf_2485,cstatus_csv_dumper_2485);
    fifo_csv_dumper_2486 = new("./depth2486.csv");
    cstatus_csv_dumper_2486 = new("./chan_status2486.csv");
    fifo_monitor_2486 = new(fifo_csv_dumper_2486,fifo_intf_2486,cstatus_csv_dumper_2486);
    fifo_csv_dumper_2487 = new("./depth2487.csv");
    cstatus_csv_dumper_2487 = new("./chan_status2487.csv");
    fifo_monitor_2487 = new(fifo_csv_dumper_2487,fifo_intf_2487,cstatus_csv_dumper_2487);
    fifo_csv_dumper_2488 = new("./depth2488.csv");
    cstatus_csv_dumper_2488 = new("./chan_status2488.csv");
    fifo_monitor_2488 = new(fifo_csv_dumper_2488,fifo_intf_2488,cstatus_csv_dumper_2488);
    fifo_csv_dumper_2489 = new("./depth2489.csv");
    cstatus_csv_dumper_2489 = new("./chan_status2489.csv");
    fifo_monitor_2489 = new(fifo_csv_dumper_2489,fifo_intf_2489,cstatus_csv_dumper_2489);
    fifo_csv_dumper_2490 = new("./depth2490.csv");
    cstatus_csv_dumper_2490 = new("./chan_status2490.csv");
    fifo_monitor_2490 = new(fifo_csv_dumper_2490,fifo_intf_2490,cstatus_csv_dumper_2490);
    fifo_csv_dumper_2491 = new("./depth2491.csv");
    cstatus_csv_dumper_2491 = new("./chan_status2491.csv");
    fifo_monitor_2491 = new(fifo_csv_dumper_2491,fifo_intf_2491,cstatus_csv_dumper_2491);
    fifo_csv_dumper_2492 = new("./depth2492.csv");
    cstatus_csv_dumper_2492 = new("./chan_status2492.csv");
    fifo_monitor_2492 = new(fifo_csv_dumper_2492,fifo_intf_2492,cstatus_csv_dumper_2492);
    fifo_csv_dumper_2493 = new("./depth2493.csv");
    cstatus_csv_dumper_2493 = new("./chan_status2493.csv");
    fifo_monitor_2493 = new(fifo_csv_dumper_2493,fifo_intf_2493,cstatus_csv_dumper_2493);
    fifo_csv_dumper_2494 = new("./depth2494.csv");
    cstatus_csv_dumper_2494 = new("./chan_status2494.csv");
    fifo_monitor_2494 = new(fifo_csv_dumper_2494,fifo_intf_2494,cstatus_csv_dumper_2494);
    fifo_csv_dumper_2495 = new("./depth2495.csv");
    cstatus_csv_dumper_2495 = new("./chan_status2495.csv");
    fifo_monitor_2495 = new(fifo_csv_dumper_2495,fifo_intf_2495,cstatus_csv_dumper_2495);
    fifo_csv_dumper_2496 = new("./depth2496.csv");
    cstatus_csv_dumper_2496 = new("./chan_status2496.csv");
    fifo_monitor_2496 = new(fifo_csv_dumper_2496,fifo_intf_2496,cstatus_csv_dumper_2496);
    fifo_csv_dumper_2497 = new("./depth2497.csv");
    cstatus_csv_dumper_2497 = new("./chan_status2497.csv");
    fifo_monitor_2497 = new(fifo_csv_dumper_2497,fifo_intf_2497,cstatus_csv_dumper_2497);
    fifo_csv_dumper_2498 = new("./depth2498.csv");
    cstatus_csv_dumper_2498 = new("./chan_status2498.csv");
    fifo_monitor_2498 = new(fifo_csv_dumper_2498,fifo_intf_2498,cstatus_csv_dumper_2498);
    fifo_csv_dumper_2499 = new("./depth2499.csv");
    cstatus_csv_dumper_2499 = new("./chan_status2499.csv");
    fifo_monitor_2499 = new(fifo_csv_dumper_2499,fifo_intf_2499,cstatus_csv_dumper_2499);
    fifo_csv_dumper_2500 = new("./depth2500.csv");
    cstatus_csv_dumper_2500 = new("./chan_status2500.csv");
    fifo_monitor_2500 = new(fifo_csv_dumper_2500,fifo_intf_2500,cstatus_csv_dumper_2500);
    fifo_csv_dumper_2501 = new("./depth2501.csv");
    cstatus_csv_dumper_2501 = new("./chan_status2501.csv");
    fifo_monitor_2501 = new(fifo_csv_dumper_2501,fifo_intf_2501,cstatus_csv_dumper_2501);
    fifo_csv_dumper_2502 = new("./depth2502.csv");
    cstatus_csv_dumper_2502 = new("./chan_status2502.csv");
    fifo_monitor_2502 = new(fifo_csv_dumper_2502,fifo_intf_2502,cstatus_csv_dumper_2502);
    fifo_csv_dumper_2503 = new("./depth2503.csv");
    cstatus_csv_dumper_2503 = new("./chan_status2503.csv");
    fifo_monitor_2503 = new(fifo_csv_dumper_2503,fifo_intf_2503,cstatus_csv_dumper_2503);
    fifo_csv_dumper_2504 = new("./depth2504.csv");
    cstatus_csv_dumper_2504 = new("./chan_status2504.csv");
    fifo_monitor_2504 = new(fifo_csv_dumper_2504,fifo_intf_2504,cstatus_csv_dumper_2504);
    fifo_csv_dumper_2505 = new("./depth2505.csv");
    cstatus_csv_dumper_2505 = new("./chan_status2505.csv");
    fifo_monitor_2505 = new(fifo_csv_dumper_2505,fifo_intf_2505,cstatus_csv_dumper_2505);
    fifo_csv_dumper_2506 = new("./depth2506.csv");
    cstatus_csv_dumper_2506 = new("./chan_status2506.csv");
    fifo_monitor_2506 = new(fifo_csv_dumper_2506,fifo_intf_2506,cstatus_csv_dumper_2506);
    fifo_csv_dumper_2507 = new("./depth2507.csv");
    cstatus_csv_dumper_2507 = new("./chan_status2507.csv");
    fifo_monitor_2507 = new(fifo_csv_dumper_2507,fifo_intf_2507,cstatus_csv_dumper_2507);
    fifo_csv_dumper_2508 = new("./depth2508.csv");
    cstatus_csv_dumper_2508 = new("./chan_status2508.csv");
    fifo_monitor_2508 = new(fifo_csv_dumper_2508,fifo_intf_2508,cstatus_csv_dumper_2508);
    fifo_csv_dumper_2509 = new("./depth2509.csv");
    cstatus_csv_dumper_2509 = new("./chan_status2509.csv");
    fifo_monitor_2509 = new(fifo_csv_dumper_2509,fifo_intf_2509,cstatus_csv_dumper_2509);
    fifo_csv_dumper_2510 = new("./depth2510.csv");
    cstatus_csv_dumper_2510 = new("./chan_status2510.csv");
    fifo_monitor_2510 = new(fifo_csv_dumper_2510,fifo_intf_2510,cstatus_csv_dumper_2510);
    fifo_csv_dumper_2511 = new("./depth2511.csv");
    cstatus_csv_dumper_2511 = new("./chan_status2511.csv");
    fifo_monitor_2511 = new(fifo_csv_dumper_2511,fifo_intf_2511,cstatus_csv_dumper_2511);
    fifo_csv_dumper_2512 = new("./depth2512.csv");
    cstatus_csv_dumper_2512 = new("./chan_status2512.csv");
    fifo_monitor_2512 = new(fifo_csv_dumper_2512,fifo_intf_2512,cstatus_csv_dumper_2512);
    fifo_csv_dumper_2513 = new("./depth2513.csv");
    cstatus_csv_dumper_2513 = new("./chan_status2513.csv");
    fifo_monitor_2513 = new(fifo_csv_dumper_2513,fifo_intf_2513,cstatus_csv_dumper_2513);
    fifo_csv_dumper_2514 = new("./depth2514.csv");
    cstatus_csv_dumper_2514 = new("./chan_status2514.csv");
    fifo_monitor_2514 = new(fifo_csv_dumper_2514,fifo_intf_2514,cstatus_csv_dumper_2514);
    fifo_csv_dumper_2515 = new("./depth2515.csv");
    cstatus_csv_dumper_2515 = new("./chan_status2515.csv");
    fifo_monitor_2515 = new(fifo_csv_dumper_2515,fifo_intf_2515,cstatus_csv_dumper_2515);
    fifo_csv_dumper_2516 = new("./depth2516.csv");
    cstatus_csv_dumper_2516 = new("./chan_status2516.csv");
    fifo_monitor_2516 = new(fifo_csv_dumper_2516,fifo_intf_2516,cstatus_csv_dumper_2516);
    fifo_csv_dumper_2517 = new("./depth2517.csv");
    cstatus_csv_dumper_2517 = new("./chan_status2517.csv");
    fifo_monitor_2517 = new(fifo_csv_dumper_2517,fifo_intf_2517,cstatus_csv_dumper_2517);
    fifo_csv_dumper_2518 = new("./depth2518.csv");
    cstatus_csv_dumper_2518 = new("./chan_status2518.csv");
    fifo_monitor_2518 = new(fifo_csv_dumper_2518,fifo_intf_2518,cstatus_csv_dumper_2518);
    fifo_csv_dumper_2519 = new("./depth2519.csv");
    cstatus_csv_dumper_2519 = new("./chan_status2519.csv");
    fifo_monitor_2519 = new(fifo_csv_dumper_2519,fifo_intf_2519,cstatus_csv_dumper_2519);
    fifo_csv_dumper_2520 = new("./depth2520.csv");
    cstatus_csv_dumper_2520 = new("./chan_status2520.csv");
    fifo_monitor_2520 = new(fifo_csv_dumper_2520,fifo_intf_2520,cstatus_csv_dumper_2520);
    fifo_csv_dumper_2521 = new("./depth2521.csv");
    cstatus_csv_dumper_2521 = new("./chan_status2521.csv");
    fifo_monitor_2521 = new(fifo_csv_dumper_2521,fifo_intf_2521,cstatus_csv_dumper_2521);
    fifo_csv_dumper_2522 = new("./depth2522.csv");
    cstatus_csv_dumper_2522 = new("./chan_status2522.csv");
    fifo_monitor_2522 = new(fifo_csv_dumper_2522,fifo_intf_2522,cstatus_csv_dumper_2522);
    fifo_csv_dumper_2523 = new("./depth2523.csv");
    cstatus_csv_dumper_2523 = new("./chan_status2523.csv");
    fifo_monitor_2523 = new(fifo_csv_dumper_2523,fifo_intf_2523,cstatus_csv_dumper_2523);
    fifo_csv_dumper_2524 = new("./depth2524.csv");
    cstatus_csv_dumper_2524 = new("./chan_status2524.csv");
    fifo_monitor_2524 = new(fifo_csv_dumper_2524,fifo_intf_2524,cstatus_csv_dumper_2524);
    fifo_csv_dumper_2525 = new("./depth2525.csv");
    cstatus_csv_dumper_2525 = new("./chan_status2525.csv");
    fifo_monitor_2525 = new(fifo_csv_dumper_2525,fifo_intf_2525,cstatus_csv_dumper_2525);
    fifo_csv_dumper_2526 = new("./depth2526.csv");
    cstatus_csv_dumper_2526 = new("./chan_status2526.csv");
    fifo_monitor_2526 = new(fifo_csv_dumper_2526,fifo_intf_2526,cstatus_csv_dumper_2526);
    fifo_csv_dumper_2527 = new("./depth2527.csv");
    cstatus_csv_dumper_2527 = new("./chan_status2527.csv");
    fifo_monitor_2527 = new(fifo_csv_dumper_2527,fifo_intf_2527,cstatus_csv_dumper_2527);
    fifo_csv_dumper_2528 = new("./depth2528.csv");
    cstatus_csv_dumper_2528 = new("./chan_status2528.csv");
    fifo_monitor_2528 = new(fifo_csv_dumper_2528,fifo_intf_2528,cstatus_csv_dumper_2528);
    fifo_csv_dumper_2529 = new("./depth2529.csv");
    cstatus_csv_dumper_2529 = new("./chan_status2529.csv");
    fifo_monitor_2529 = new(fifo_csv_dumper_2529,fifo_intf_2529,cstatus_csv_dumper_2529);
    fifo_csv_dumper_2530 = new("./depth2530.csv");
    cstatus_csv_dumper_2530 = new("./chan_status2530.csv");
    fifo_monitor_2530 = new(fifo_csv_dumper_2530,fifo_intf_2530,cstatus_csv_dumper_2530);
    fifo_csv_dumper_2531 = new("./depth2531.csv");
    cstatus_csv_dumper_2531 = new("./chan_status2531.csv");
    fifo_monitor_2531 = new(fifo_csv_dumper_2531,fifo_intf_2531,cstatus_csv_dumper_2531);
    fifo_csv_dumper_2532 = new("./depth2532.csv");
    cstatus_csv_dumper_2532 = new("./chan_status2532.csv");
    fifo_monitor_2532 = new(fifo_csv_dumper_2532,fifo_intf_2532,cstatus_csv_dumper_2532);
    fifo_csv_dumper_2533 = new("./depth2533.csv");
    cstatus_csv_dumper_2533 = new("./chan_status2533.csv");
    fifo_monitor_2533 = new(fifo_csv_dumper_2533,fifo_intf_2533,cstatus_csv_dumper_2533);
    fifo_csv_dumper_2534 = new("./depth2534.csv");
    cstatus_csv_dumper_2534 = new("./chan_status2534.csv");
    fifo_monitor_2534 = new(fifo_csv_dumper_2534,fifo_intf_2534,cstatus_csv_dumper_2534);
    fifo_csv_dumper_2535 = new("./depth2535.csv");
    cstatus_csv_dumper_2535 = new("./chan_status2535.csv");
    fifo_monitor_2535 = new(fifo_csv_dumper_2535,fifo_intf_2535,cstatus_csv_dumper_2535);
    fifo_csv_dumper_2536 = new("./depth2536.csv");
    cstatus_csv_dumper_2536 = new("./chan_status2536.csv");
    fifo_monitor_2536 = new(fifo_csv_dumper_2536,fifo_intf_2536,cstatus_csv_dumper_2536);
    fifo_csv_dumper_2537 = new("./depth2537.csv");
    cstatus_csv_dumper_2537 = new("./chan_status2537.csv");
    fifo_monitor_2537 = new(fifo_csv_dumper_2537,fifo_intf_2537,cstatus_csv_dumper_2537);
    fifo_csv_dumper_2538 = new("./depth2538.csv");
    cstatus_csv_dumper_2538 = new("./chan_status2538.csv");
    fifo_monitor_2538 = new(fifo_csv_dumper_2538,fifo_intf_2538,cstatus_csv_dumper_2538);
    fifo_csv_dumper_2539 = new("./depth2539.csv");
    cstatus_csv_dumper_2539 = new("./chan_status2539.csv");
    fifo_monitor_2539 = new(fifo_csv_dumper_2539,fifo_intf_2539,cstatus_csv_dumper_2539);
    fifo_csv_dumper_2540 = new("./depth2540.csv");
    cstatus_csv_dumper_2540 = new("./chan_status2540.csv");
    fifo_monitor_2540 = new(fifo_csv_dumper_2540,fifo_intf_2540,cstatus_csv_dumper_2540);
    fifo_csv_dumper_2541 = new("./depth2541.csv");
    cstatus_csv_dumper_2541 = new("./chan_status2541.csv");
    fifo_monitor_2541 = new(fifo_csv_dumper_2541,fifo_intf_2541,cstatus_csv_dumper_2541);
    fifo_csv_dumper_2542 = new("./depth2542.csv");
    cstatus_csv_dumper_2542 = new("./chan_status2542.csv");
    fifo_monitor_2542 = new(fifo_csv_dumper_2542,fifo_intf_2542,cstatus_csv_dumper_2542);
    fifo_csv_dumper_2543 = new("./depth2543.csv");
    cstatus_csv_dumper_2543 = new("./chan_status2543.csv");
    fifo_monitor_2543 = new(fifo_csv_dumper_2543,fifo_intf_2543,cstatus_csv_dumper_2543);
    fifo_csv_dumper_2544 = new("./depth2544.csv");
    cstatus_csv_dumper_2544 = new("./chan_status2544.csv");
    fifo_monitor_2544 = new(fifo_csv_dumper_2544,fifo_intf_2544,cstatus_csv_dumper_2544);
    fifo_csv_dumper_2545 = new("./depth2545.csv");
    cstatus_csv_dumper_2545 = new("./chan_status2545.csv");
    fifo_monitor_2545 = new(fifo_csv_dumper_2545,fifo_intf_2545,cstatus_csv_dumper_2545);
    fifo_csv_dumper_2546 = new("./depth2546.csv");
    cstatus_csv_dumper_2546 = new("./chan_status2546.csv");
    fifo_monitor_2546 = new(fifo_csv_dumper_2546,fifo_intf_2546,cstatus_csv_dumper_2546);
    fifo_csv_dumper_2547 = new("./depth2547.csv");
    cstatus_csv_dumper_2547 = new("./chan_status2547.csv");
    fifo_monitor_2547 = new(fifo_csv_dumper_2547,fifo_intf_2547,cstatus_csv_dumper_2547);
    fifo_csv_dumper_2548 = new("./depth2548.csv");
    cstatus_csv_dumper_2548 = new("./chan_status2548.csv");
    fifo_monitor_2548 = new(fifo_csv_dumper_2548,fifo_intf_2548,cstatus_csv_dumper_2548);
    fifo_csv_dumper_2549 = new("./depth2549.csv");
    cstatus_csv_dumper_2549 = new("./chan_status2549.csv");
    fifo_monitor_2549 = new(fifo_csv_dumper_2549,fifo_intf_2549,cstatus_csv_dumper_2549);
    fifo_csv_dumper_2550 = new("./depth2550.csv");
    cstatus_csv_dumper_2550 = new("./chan_status2550.csv");
    fifo_monitor_2550 = new(fifo_csv_dumper_2550,fifo_intf_2550,cstatus_csv_dumper_2550);
    fifo_csv_dumper_2551 = new("./depth2551.csv");
    cstatus_csv_dumper_2551 = new("./chan_status2551.csv");
    fifo_monitor_2551 = new(fifo_csv_dumper_2551,fifo_intf_2551,cstatus_csv_dumper_2551);
    fifo_csv_dumper_2552 = new("./depth2552.csv");
    cstatus_csv_dumper_2552 = new("./chan_status2552.csv");
    fifo_monitor_2552 = new(fifo_csv_dumper_2552,fifo_intf_2552,cstatus_csv_dumper_2552);
    fifo_csv_dumper_2553 = new("./depth2553.csv");
    cstatus_csv_dumper_2553 = new("./chan_status2553.csv");
    fifo_monitor_2553 = new(fifo_csv_dumper_2553,fifo_intf_2553,cstatus_csv_dumper_2553);
    fifo_csv_dumper_2554 = new("./depth2554.csv");
    cstatus_csv_dumper_2554 = new("./chan_status2554.csv");
    fifo_monitor_2554 = new(fifo_csv_dumper_2554,fifo_intf_2554,cstatus_csv_dumper_2554);
    fifo_csv_dumper_2555 = new("./depth2555.csv");
    cstatus_csv_dumper_2555 = new("./chan_status2555.csv");
    fifo_monitor_2555 = new(fifo_csv_dumper_2555,fifo_intf_2555,cstatus_csv_dumper_2555);
    fifo_csv_dumper_2556 = new("./depth2556.csv");
    cstatus_csv_dumper_2556 = new("./chan_status2556.csv");
    fifo_monitor_2556 = new(fifo_csv_dumper_2556,fifo_intf_2556,cstatus_csv_dumper_2556);
    fifo_csv_dumper_2557 = new("./depth2557.csv");
    cstatus_csv_dumper_2557 = new("./chan_status2557.csv");
    fifo_monitor_2557 = new(fifo_csv_dumper_2557,fifo_intf_2557,cstatus_csv_dumper_2557);
    fifo_csv_dumper_2558 = new("./depth2558.csv");
    cstatus_csv_dumper_2558 = new("./chan_status2558.csv");
    fifo_monitor_2558 = new(fifo_csv_dumper_2558,fifo_intf_2558,cstatus_csv_dumper_2558);
    fifo_csv_dumper_2559 = new("./depth2559.csv");
    cstatus_csv_dumper_2559 = new("./chan_status2559.csv");
    fifo_monitor_2559 = new(fifo_csv_dumper_2559,fifo_intf_2559,cstatus_csv_dumper_2559);
    fifo_csv_dumper_2560 = new("./depth2560.csv");
    cstatus_csv_dumper_2560 = new("./chan_status2560.csv");
    fifo_monitor_2560 = new(fifo_csv_dumper_2560,fifo_intf_2560,cstatus_csv_dumper_2560);
    fifo_csv_dumper_2561 = new("./depth2561.csv");
    cstatus_csv_dumper_2561 = new("./chan_status2561.csv");
    fifo_monitor_2561 = new(fifo_csv_dumper_2561,fifo_intf_2561,cstatus_csv_dumper_2561);
    fifo_csv_dumper_2562 = new("./depth2562.csv");
    cstatus_csv_dumper_2562 = new("./chan_status2562.csv");
    fifo_monitor_2562 = new(fifo_csv_dumper_2562,fifo_intf_2562,cstatus_csv_dumper_2562);
    fifo_csv_dumper_2563 = new("./depth2563.csv");
    cstatus_csv_dumper_2563 = new("./chan_status2563.csv");
    fifo_monitor_2563 = new(fifo_csv_dumper_2563,fifo_intf_2563,cstatus_csv_dumper_2563);
    fifo_csv_dumper_2564 = new("./depth2564.csv");
    cstatus_csv_dumper_2564 = new("./chan_status2564.csv");
    fifo_monitor_2564 = new(fifo_csv_dumper_2564,fifo_intf_2564,cstatus_csv_dumper_2564);
    fifo_csv_dumper_2565 = new("./depth2565.csv");
    cstatus_csv_dumper_2565 = new("./chan_status2565.csv");
    fifo_monitor_2565 = new(fifo_csv_dumper_2565,fifo_intf_2565,cstatus_csv_dumper_2565);
    fifo_csv_dumper_2566 = new("./depth2566.csv");
    cstatus_csv_dumper_2566 = new("./chan_status2566.csv");
    fifo_monitor_2566 = new(fifo_csv_dumper_2566,fifo_intf_2566,cstatus_csv_dumper_2566);
    fifo_csv_dumper_2567 = new("./depth2567.csv");
    cstatus_csv_dumper_2567 = new("./chan_status2567.csv");
    fifo_monitor_2567 = new(fifo_csv_dumper_2567,fifo_intf_2567,cstatus_csv_dumper_2567);
    fifo_csv_dumper_2568 = new("./depth2568.csv");
    cstatus_csv_dumper_2568 = new("./chan_status2568.csv");
    fifo_monitor_2568 = new(fifo_csv_dumper_2568,fifo_intf_2568,cstatus_csv_dumper_2568);
    fifo_csv_dumper_2569 = new("./depth2569.csv");
    cstatus_csv_dumper_2569 = new("./chan_status2569.csv");
    fifo_monitor_2569 = new(fifo_csv_dumper_2569,fifo_intf_2569,cstatus_csv_dumper_2569);
    fifo_csv_dumper_2570 = new("./depth2570.csv");
    cstatus_csv_dumper_2570 = new("./chan_status2570.csv");
    fifo_monitor_2570 = new(fifo_csv_dumper_2570,fifo_intf_2570,cstatus_csv_dumper_2570);
    fifo_csv_dumper_2571 = new("./depth2571.csv");
    cstatus_csv_dumper_2571 = new("./chan_status2571.csv");
    fifo_monitor_2571 = new(fifo_csv_dumper_2571,fifo_intf_2571,cstatus_csv_dumper_2571);
    fifo_csv_dumper_2572 = new("./depth2572.csv");
    cstatus_csv_dumper_2572 = new("./chan_status2572.csv");
    fifo_monitor_2572 = new(fifo_csv_dumper_2572,fifo_intf_2572,cstatus_csv_dumper_2572);
    fifo_csv_dumper_2573 = new("./depth2573.csv");
    cstatus_csv_dumper_2573 = new("./chan_status2573.csv");
    fifo_monitor_2573 = new(fifo_csv_dumper_2573,fifo_intf_2573,cstatus_csv_dumper_2573);
    fifo_csv_dumper_2574 = new("./depth2574.csv");
    cstatus_csv_dumper_2574 = new("./chan_status2574.csv");
    fifo_monitor_2574 = new(fifo_csv_dumper_2574,fifo_intf_2574,cstatus_csv_dumper_2574);
    fifo_csv_dumper_2575 = new("./depth2575.csv");
    cstatus_csv_dumper_2575 = new("./chan_status2575.csv");
    fifo_monitor_2575 = new(fifo_csv_dumper_2575,fifo_intf_2575,cstatus_csv_dumper_2575);
    fifo_csv_dumper_2576 = new("./depth2576.csv");
    cstatus_csv_dumper_2576 = new("./chan_status2576.csv");
    fifo_monitor_2576 = new(fifo_csv_dumper_2576,fifo_intf_2576,cstatus_csv_dumper_2576);
    fifo_csv_dumper_2577 = new("./depth2577.csv");
    cstatus_csv_dumper_2577 = new("./chan_status2577.csv");
    fifo_monitor_2577 = new(fifo_csv_dumper_2577,fifo_intf_2577,cstatus_csv_dumper_2577);
    fifo_csv_dumper_2578 = new("./depth2578.csv");
    cstatus_csv_dumper_2578 = new("./chan_status2578.csv");
    fifo_monitor_2578 = new(fifo_csv_dumper_2578,fifo_intf_2578,cstatus_csv_dumper_2578);
    fifo_csv_dumper_2579 = new("./depth2579.csv");
    cstatus_csv_dumper_2579 = new("./chan_status2579.csv");
    fifo_monitor_2579 = new(fifo_csv_dumper_2579,fifo_intf_2579,cstatus_csv_dumper_2579);
    fifo_csv_dumper_2580 = new("./depth2580.csv");
    cstatus_csv_dumper_2580 = new("./chan_status2580.csv");
    fifo_monitor_2580 = new(fifo_csv_dumper_2580,fifo_intf_2580,cstatus_csv_dumper_2580);
    fifo_csv_dumper_2581 = new("./depth2581.csv");
    cstatus_csv_dumper_2581 = new("./chan_status2581.csv");
    fifo_monitor_2581 = new(fifo_csv_dumper_2581,fifo_intf_2581,cstatus_csv_dumper_2581);
    fifo_csv_dumper_2582 = new("./depth2582.csv");
    cstatus_csv_dumper_2582 = new("./chan_status2582.csv");
    fifo_monitor_2582 = new(fifo_csv_dumper_2582,fifo_intf_2582,cstatus_csv_dumper_2582);
    fifo_csv_dumper_2583 = new("./depth2583.csv");
    cstatus_csv_dumper_2583 = new("./chan_status2583.csv");
    fifo_monitor_2583 = new(fifo_csv_dumper_2583,fifo_intf_2583,cstatus_csv_dumper_2583);
    fifo_csv_dumper_2584 = new("./depth2584.csv");
    cstatus_csv_dumper_2584 = new("./chan_status2584.csv");
    fifo_monitor_2584 = new(fifo_csv_dumper_2584,fifo_intf_2584,cstatus_csv_dumper_2584);
    fifo_csv_dumper_2585 = new("./depth2585.csv");
    cstatus_csv_dumper_2585 = new("./chan_status2585.csv");
    fifo_monitor_2585 = new(fifo_csv_dumper_2585,fifo_intf_2585,cstatus_csv_dumper_2585);
    fifo_csv_dumper_2586 = new("./depth2586.csv");
    cstatus_csv_dumper_2586 = new("./chan_status2586.csv");
    fifo_monitor_2586 = new(fifo_csv_dumper_2586,fifo_intf_2586,cstatus_csv_dumper_2586);
    fifo_csv_dumper_2587 = new("./depth2587.csv");
    cstatus_csv_dumper_2587 = new("./chan_status2587.csv");
    fifo_monitor_2587 = new(fifo_csv_dumper_2587,fifo_intf_2587,cstatus_csv_dumper_2587);
    fifo_csv_dumper_2588 = new("./depth2588.csv");
    cstatus_csv_dumper_2588 = new("./chan_status2588.csv");
    fifo_monitor_2588 = new(fifo_csv_dumper_2588,fifo_intf_2588,cstatus_csv_dumper_2588);
    fifo_csv_dumper_2589 = new("./depth2589.csv");
    cstatus_csv_dumper_2589 = new("./chan_status2589.csv");
    fifo_monitor_2589 = new(fifo_csv_dumper_2589,fifo_intf_2589,cstatus_csv_dumper_2589);
    fifo_csv_dumper_2590 = new("./depth2590.csv");
    cstatus_csv_dumper_2590 = new("./chan_status2590.csv");
    fifo_monitor_2590 = new(fifo_csv_dumper_2590,fifo_intf_2590,cstatus_csv_dumper_2590);
    fifo_csv_dumper_2591 = new("./depth2591.csv");
    cstatus_csv_dumper_2591 = new("./chan_status2591.csv");
    fifo_monitor_2591 = new(fifo_csv_dumper_2591,fifo_intf_2591,cstatus_csv_dumper_2591);
    fifo_csv_dumper_2592 = new("./depth2592.csv");
    cstatus_csv_dumper_2592 = new("./chan_status2592.csv");
    fifo_monitor_2592 = new(fifo_csv_dumper_2592,fifo_intf_2592,cstatus_csv_dumper_2592);
    fifo_csv_dumper_2593 = new("./depth2593.csv");
    cstatus_csv_dumper_2593 = new("./chan_status2593.csv");
    fifo_monitor_2593 = new(fifo_csv_dumper_2593,fifo_intf_2593,cstatus_csv_dumper_2593);
    fifo_csv_dumper_2594 = new("./depth2594.csv");
    cstatus_csv_dumper_2594 = new("./chan_status2594.csv");
    fifo_monitor_2594 = new(fifo_csv_dumper_2594,fifo_intf_2594,cstatus_csv_dumper_2594);
    fifo_csv_dumper_2595 = new("./depth2595.csv");
    cstatus_csv_dumper_2595 = new("./chan_status2595.csv");
    fifo_monitor_2595 = new(fifo_csv_dumper_2595,fifo_intf_2595,cstatus_csv_dumper_2595);
    fifo_csv_dumper_2596 = new("./depth2596.csv");
    cstatus_csv_dumper_2596 = new("./chan_status2596.csv");
    fifo_monitor_2596 = new(fifo_csv_dumper_2596,fifo_intf_2596,cstatus_csv_dumper_2596);
    fifo_csv_dumper_2597 = new("./depth2597.csv");
    cstatus_csv_dumper_2597 = new("./chan_status2597.csv");
    fifo_monitor_2597 = new(fifo_csv_dumper_2597,fifo_intf_2597,cstatus_csv_dumper_2597);
    fifo_csv_dumper_2598 = new("./depth2598.csv");
    cstatus_csv_dumper_2598 = new("./chan_status2598.csv");
    fifo_monitor_2598 = new(fifo_csv_dumper_2598,fifo_intf_2598,cstatus_csv_dumper_2598);
    fifo_csv_dumper_2599 = new("./depth2599.csv");
    cstatus_csv_dumper_2599 = new("./chan_status2599.csv");
    fifo_monitor_2599 = new(fifo_csv_dumper_2599,fifo_intf_2599,cstatus_csv_dumper_2599);
    fifo_csv_dumper_2600 = new("./depth2600.csv");
    cstatus_csv_dumper_2600 = new("./chan_status2600.csv");
    fifo_monitor_2600 = new(fifo_csv_dumper_2600,fifo_intf_2600,cstatus_csv_dumper_2600);
    fifo_csv_dumper_2601 = new("./depth2601.csv");
    cstatus_csv_dumper_2601 = new("./chan_status2601.csv");
    fifo_monitor_2601 = new(fifo_csv_dumper_2601,fifo_intf_2601,cstatus_csv_dumper_2601);
    fifo_csv_dumper_2602 = new("./depth2602.csv");
    cstatus_csv_dumper_2602 = new("./chan_status2602.csv");
    fifo_monitor_2602 = new(fifo_csv_dumper_2602,fifo_intf_2602,cstatus_csv_dumper_2602);
    fifo_csv_dumper_2603 = new("./depth2603.csv");
    cstatus_csv_dumper_2603 = new("./chan_status2603.csv");
    fifo_monitor_2603 = new(fifo_csv_dumper_2603,fifo_intf_2603,cstatus_csv_dumper_2603);
    fifo_csv_dumper_2604 = new("./depth2604.csv");
    cstatus_csv_dumper_2604 = new("./chan_status2604.csv");
    fifo_monitor_2604 = new(fifo_csv_dumper_2604,fifo_intf_2604,cstatus_csv_dumper_2604);
    fifo_csv_dumper_2605 = new("./depth2605.csv");
    cstatus_csv_dumper_2605 = new("./chan_status2605.csv");
    fifo_monitor_2605 = new(fifo_csv_dumper_2605,fifo_intf_2605,cstatus_csv_dumper_2605);
    fifo_csv_dumper_2606 = new("./depth2606.csv");
    cstatus_csv_dumper_2606 = new("./chan_status2606.csv");
    fifo_monitor_2606 = new(fifo_csv_dumper_2606,fifo_intf_2606,cstatus_csv_dumper_2606);
    fifo_csv_dumper_2607 = new("./depth2607.csv");
    cstatus_csv_dumper_2607 = new("./chan_status2607.csv");
    fifo_monitor_2607 = new(fifo_csv_dumper_2607,fifo_intf_2607,cstatus_csv_dumper_2607);
    fifo_csv_dumper_2608 = new("./depth2608.csv");
    cstatus_csv_dumper_2608 = new("./chan_status2608.csv");
    fifo_monitor_2608 = new(fifo_csv_dumper_2608,fifo_intf_2608,cstatus_csv_dumper_2608);
    fifo_csv_dumper_2609 = new("./depth2609.csv");
    cstatus_csv_dumper_2609 = new("./chan_status2609.csv");
    fifo_monitor_2609 = new(fifo_csv_dumper_2609,fifo_intf_2609,cstatus_csv_dumper_2609);
    fifo_csv_dumper_2610 = new("./depth2610.csv");
    cstatus_csv_dumper_2610 = new("./chan_status2610.csv");
    fifo_monitor_2610 = new(fifo_csv_dumper_2610,fifo_intf_2610,cstatus_csv_dumper_2610);
    fifo_csv_dumper_2611 = new("./depth2611.csv");
    cstatus_csv_dumper_2611 = new("./chan_status2611.csv");
    fifo_monitor_2611 = new(fifo_csv_dumper_2611,fifo_intf_2611,cstatus_csv_dumper_2611);
    fifo_csv_dumper_2612 = new("./depth2612.csv");
    cstatus_csv_dumper_2612 = new("./chan_status2612.csv");
    fifo_monitor_2612 = new(fifo_csv_dumper_2612,fifo_intf_2612,cstatus_csv_dumper_2612);
    fifo_csv_dumper_2613 = new("./depth2613.csv");
    cstatus_csv_dumper_2613 = new("./chan_status2613.csv");
    fifo_monitor_2613 = new(fifo_csv_dumper_2613,fifo_intf_2613,cstatus_csv_dumper_2613);
    fifo_csv_dumper_2614 = new("./depth2614.csv");
    cstatus_csv_dumper_2614 = new("./chan_status2614.csv");
    fifo_monitor_2614 = new(fifo_csv_dumper_2614,fifo_intf_2614,cstatus_csv_dumper_2614);
    fifo_csv_dumper_2615 = new("./depth2615.csv");
    cstatus_csv_dumper_2615 = new("./chan_status2615.csv");
    fifo_monitor_2615 = new(fifo_csv_dumper_2615,fifo_intf_2615,cstatus_csv_dumper_2615);
    fifo_csv_dumper_2616 = new("./depth2616.csv");
    cstatus_csv_dumper_2616 = new("./chan_status2616.csv");
    fifo_monitor_2616 = new(fifo_csv_dumper_2616,fifo_intf_2616,cstatus_csv_dumper_2616);
    fifo_csv_dumper_2617 = new("./depth2617.csv");
    cstatus_csv_dumper_2617 = new("./chan_status2617.csv");
    fifo_monitor_2617 = new(fifo_csv_dumper_2617,fifo_intf_2617,cstatus_csv_dumper_2617);
    fifo_csv_dumper_2618 = new("./depth2618.csv");
    cstatus_csv_dumper_2618 = new("./chan_status2618.csv");
    fifo_monitor_2618 = new(fifo_csv_dumper_2618,fifo_intf_2618,cstatus_csv_dumper_2618);
    fifo_csv_dumper_2619 = new("./depth2619.csv");
    cstatus_csv_dumper_2619 = new("./chan_status2619.csv");
    fifo_monitor_2619 = new(fifo_csv_dumper_2619,fifo_intf_2619,cstatus_csv_dumper_2619);
    fifo_csv_dumper_2620 = new("./depth2620.csv");
    cstatus_csv_dumper_2620 = new("./chan_status2620.csv");
    fifo_monitor_2620 = new(fifo_csv_dumper_2620,fifo_intf_2620,cstatus_csv_dumper_2620);
    fifo_csv_dumper_2621 = new("./depth2621.csv");
    cstatus_csv_dumper_2621 = new("./chan_status2621.csv");
    fifo_monitor_2621 = new(fifo_csv_dumper_2621,fifo_intf_2621,cstatus_csv_dumper_2621);
    fifo_csv_dumper_2622 = new("./depth2622.csv");
    cstatus_csv_dumper_2622 = new("./chan_status2622.csv");
    fifo_monitor_2622 = new(fifo_csv_dumper_2622,fifo_intf_2622,cstatus_csv_dumper_2622);
    fifo_csv_dumper_2623 = new("./depth2623.csv");
    cstatus_csv_dumper_2623 = new("./chan_status2623.csv");
    fifo_monitor_2623 = new(fifo_csv_dumper_2623,fifo_intf_2623,cstatus_csv_dumper_2623);
    fifo_csv_dumper_2624 = new("./depth2624.csv");
    cstatus_csv_dumper_2624 = new("./chan_status2624.csv");
    fifo_monitor_2624 = new(fifo_csv_dumper_2624,fifo_intf_2624,cstatus_csv_dumper_2624);
    fifo_csv_dumper_2625 = new("./depth2625.csv");
    cstatus_csv_dumper_2625 = new("./chan_status2625.csv");
    fifo_monitor_2625 = new(fifo_csv_dumper_2625,fifo_intf_2625,cstatus_csv_dumper_2625);
    fifo_csv_dumper_2626 = new("./depth2626.csv");
    cstatus_csv_dumper_2626 = new("./chan_status2626.csv");
    fifo_monitor_2626 = new(fifo_csv_dumper_2626,fifo_intf_2626,cstatus_csv_dumper_2626);
    fifo_csv_dumper_2627 = new("./depth2627.csv");
    cstatus_csv_dumper_2627 = new("./chan_status2627.csv");
    fifo_monitor_2627 = new(fifo_csv_dumper_2627,fifo_intf_2627,cstatus_csv_dumper_2627);
    fifo_csv_dumper_2628 = new("./depth2628.csv");
    cstatus_csv_dumper_2628 = new("./chan_status2628.csv");
    fifo_monitor_2628 = new(fifo_csv_dumper_2628,fifo_intf_2628,cstatus_csv_dumper_2628);
    fifo_csv_dumper_2629 = new("./depth2629.csv");
    cstatus_csv_dumper_2629 = new("./chan_status2629.csv");
    fifo_monitor_2629 = new(fifo_csv_dumper_2629,fifo_intf_2629,cstatus_csv_dumper_2629);
    fifo_csv_dumper_2630 = new("./depth2630.csv");
    cstatus_csv_dumper_2630 = new("./chan_status2630.csv");
    fifo_monitor_2630 = new(fifo_csv_dumper_2630,fifo_intf_2630,cstatus_csv_dumper_2630);
    fifo_csv_dumper_2631 = new("./depth2631.csv");
    cstatus_csv_dumper_2631 = new("./chan_status2631.csv");
    fifo_monitor_2631 = new(fifo_csv_dumper_2631,fifo_intf_2631,cstatus_csv_dumper_2631);
    fifo_csv_dumper_2632 = new("./depth2632.csv");
    cstatus_csv_dumper_2632 = new("./chan_status2632.csv");
    fifo_monitor_2632 = new(fifo_csv_dumper_2632,fifo_intf_2632,cstatus_csv_dumper_2632);
    fifo_csv_dumper_2633 = new("./depth2633.csv");
    cstatus_csv_dumper_2633 = new("./chan_status2633.csv");
    fifo_monitor_2633 = new(fifo_csv_dumper_2633,fifo_intf_2633,cstatus_csv_dumper_2633);
    fifo_csv_dumper_2634 = new("./depth2634.csv");
    cstatus_csv_dumper_2634 = new("./chan_status2634.csv");
    fifo_monitor_2634 = new(fifo_csv_dumper_2634,fifo_intf_2634,cstatus_csv_dumper_2634);
    fifo_csv_dumper_2635 = new("./depth2635.csv");
    cstatus_csv_dumper_2635 = new("./chan_status2635.csv");
    fifo_monitor_2635 = new(fifo_csv_dumper_2635,fifo_intf_2635,cstatus_csv_dumper_2635);
    fifo_csv_dumper_2636 = new("./depth2636.csv");
    cstatus_csv_dumper_2636 = new("./chan_status2636.csv");
    fifo_monitor_2636 = new(fifo_csv_dumper_2636,fifo_intf_2636,cstatus_csv_dumper_2636);
    fifo_csv_dumper_2637 = new("./depth2637.csv");
    cstatus_csv_dumper_2637 = new("./chan_status2637.csv");
    fifo_monitor_2637 = new(fifo_csv_dumper_2637,fifo_intf_2637,cstatus_csv_dumper_2637);
    fifo_csv_dumper_2638 = new("./depth2638.csv");
    cstatus_csv_dumper_2638 = new("./chan_status2638.csv");
    fifo_monitor_2638 = new(fifo_csv_dumper_2638,fifo_intf_2638,cstatus_csv_dumper_2638);
    fifo_csv_dumper_2639 = new("./depth2639.csv");
    cstatus_csv_dumper_2639 = new("./chan_status2639.csv");
    fifo_monitor_2639 = new(fifo_csv_dumper_2639,fifo_intf_2639,cstatus_csv_dumper_2639);
    fifo_csv_dumper_2640 = new("./depth2640.csv");
    cstatus_csv_dumper_2640 = new("./chan_status2640.csv");
    fifo_monitor_2640 = new(fifo_csv_dumper_2640,fifo_intf_2640,cstatus_csv_dumper_2640);
    fifo_csv_dumper_2641 = new("./depth2641.csv");
    cstatus_csv_dumper_2641 = new("./chan_status2641.csv");
    fifo_monitor_2641 = new(fifo_csv_dumper_2641,fifo_intf_2641,cstatus_csv_dumper_2641);
    fifo_csv_dumper_2642 = new("./depth2642.csv");
    cstatus_csv_dumper_2642 = new("./chan_status2642.csv");
    fifo_monitor_2642 = new(fifo_csv_dumper_2642,fifo_intf_2642,cstatus_csv_dumper_2642);
    fifo_csv_dumper_2643 = new("./depth2643.csv");
    cstatus_csv_dumper_2643 = new("./chan_status2643.csv");
    fifo_monitor_2643 = new(fifo_csv_dumper_2643,fifo_intf_2643,cstatus_csv_dumper_2643);
    fifo_csv_dumper_2644 = new("./depth2644.csv");
    cstatus_csv_dumper_2644 = new("./chan_status2644.csv");
    fifo_monitor_2644 = new(fifo_csv_dumper_2644,fifo_intf_2644,cstatus_csv_dumper_2644);
    fifo_csv_dumper_2645 = new("./depth2645.csv");
    cstatus_csv_dumper_2645 = new("./chan_status2645.csv");
    fifo_monitor_2645 = new(fifo_csv_dumper_2645,fifo_intf_2645,cstatus_csv_dumper_2645);
    fifo_csv_dumper_2646 = new("./depth2646.csv");
    cstatus_csv_dumper_2646 = new("./chan_status2646.csv");
    fifo_monitor_2646 = new(fifo_csv_dumper_2646,fifo_intf_2646,cstatus_csv_dumper_2646);
    fifo_csv_dumper_2647 = new("./depth2647.csv");
    cstatus_csv_dumper_2647 = new("./chan_status2647.csv");
    fifo_monitor_2647 = new(fifo_csv_dumper_2647,fifo_intf_2647,cstatus_csv_dumper_2647);
    fifo_csv_dumper_2648 = new("./depth2648.csv");
    cstatus_csv_dumper_2648 = new("./chan_status2648.csv");
    fifo_monitor_2648 = new(fifo_csv_dumper_2648,fifo_intf_2648,cstatus_csv_dumper_2648);
    fifo_csv_dumper_2649 = new("./depth2649.csv");
    cstatus_csv_dumper_2649 = new("./chan_status2649.csv");
    fifo_monitor_2649 = new(fifo_csv_dumper_2649,fifo_intf_2649,cstatus_csv_dumper_2649);
    fifo_csv_dumper_2650 = new("./depth2650.csv");
    cstatus_csv_dumper_2650 = new("./chan_status2650.csv");
    fifo_monitor_2650 = new(fifo_csv_dumper_2650,fifo_intf_2650,cstatus_csv_dumper_2650);
    fifo_csv_dumper_2651 = new("./depth2651.csv");
    cstatus_csv_dumper_2651 = new("./chan_status2651.csv");
    fifo_monitor_2651 = new(fifo_csv_dumper_2651,fifo_intf_2651,cstatus_csv_dumper_2651);
    fifo_csv_dumper_2652 = new("./depth2652.csv");
    cstatus_csv_dumper_2652 = new("./chan_status2652.csv");
    fifo_monitor_2652 = new(fifo_csv_dumper_2652,fifo_intf_2652,cstatus_csv_dumper_2652);
    fifo_csv_dumper_2653 = new("./depth2653.csv");
    cstatus_csv_dumper_2653 = new("./chan_status2653.csv");
    fifo_monitor_2653 = new(fifo_csv_dumper_2653,fifo_intf_2653,cstatus_csv_dumper_2653);
    fifo_csv_dumper_2654 = new("./depth2654.csv");
    cstatus_csv_dumper_2654 = new("./chan_status2654.csv");
    fifo_monitor_2654 = new(fifo_csv_dumper_2654,fifo_intf_2654,cstatus_csv_dumper_2654);
    fifo_csv_dumper_2655 = new("./depth2655.csv");
    cstatus_csv_dumper_2655 = new("./chan_status2655.csv");
    fifo_monitor_2655 = new(fifo_csv_dumper_2655,fifo_intf_2655,cstatus_csv_dumper_2655);
    fifo_csv_dumper_2656 = new("./depth2656.csv");
    cstatus_csv_dumper_2656 = new("./chan_status2656.csv");
    fifo_monitor_2656 = new(fifo_csv_dumper_2656,fifo_intf_2656,cstatus_csv_dumper_2656);
    fifo_csv_dumper_2657 = new("./depth2657.csv");
    cstatus_csv_dumper_2657 = new("./chan_status2657.csv");
    fifo_monitor_2657 = new(fifo_csv_dumper_2657,fifo_intf_2657,cstatus_csv_dumper_2657);
    fifo_csv_dumper_2658 = new("./depth2658.csv");
    cstatus_csv_dumper_2658 = new("./chan_status2658.csv");
    fifo_monitor_2658 = new(fifo_csv_dumper_2658,fifo_intf_2658,cstatus_csv_dumper_2658);
    fifo_csv_dumper_2659 = new("./depth2659.csv");
    cstatus_csv_dumper_2659 = new("./chan_status2659.csv");
    fifo_monitor_2659 = new(fifo_csv_dumper_2659,fifo_intf_2659,cstatus_csv_dumper_2659);
    fifo_csv_dumper_2660 = new("./depth2660.csv");
    cstatus_csv_dumper_2660 = new("./chan_status2660.csv");
    fifo_monitor_2660 = new(fifo_csv_dumper_2660,fifo_intf_2660,cstatus_csv_dumper_2660);
    fifo_csv_dumper_2661 = new("./depth2661.csv");
    cstatus_csv_dumper_2661 = new("./chan_status2661.csv");
    fifo_monitor_2661 = new(fifo_csv_dumper_2661,fifo_intf_2661,cstatus_csv_dumper_2661);
    fifo_csv_dumper_2662 = new("./depth2662.csv");
    cstatus_csv_dumper_2662 = new("./chan_status2662.csv");
    fifo_monitor_2662 = new(fifo_csv_dumper_2662,fifo_intf_2662,cstatus_csv_dumper_2662);
    fifo_csv_dumper_2663 = new("./depth2663.csv");
    cstatus_csv_dumper_2663 = new("./chan_status2663.csv");
    fifo_monitor_2663 = new(fifo_csv_dumper_2663,fifo_intf_2663,cstatus_csv_dumper_2663);
    fifo_csv_dumper_2664 = new("./depth2664.csv");
    cstatus_csv_dumper_2664 = new("./chan_status2664.csv");
    fifo_monitor_2664 = new(fifo_csv_dumper_2664,fifo_intf_2664,cstatus_csv_dumper_2664);
    fifo_csv_dumper_2665 = new("./depth2665.csv");
    cstatus_csv_dumper_2665 = new("./chan_status2665.csv");
    fifo_monitor_2665 = new(fifo_csv_dumper_2665,fifo_intf_2665,cstatus_csv_dumper_2665);
    fifo_csv_dumper_2666 = new("./depth2666.csv");
    cstatus_csv_dumper_2666 = new("./chan_status2666.csv");
    fifo_monitor_2666 = new(fifo_csv_dumper_2666,fifo_intf_2666,cstatus_csv_dumper_2666);
    fifo_csv_dumper_2667 = new("./depth2667.csv");
    cstatus_csv_dumper_2667 = new("./chan_status2667.csv");
    fifo_monitor_2667 = new(fifo_csv_dumper_2667,fifo_intf_2667,cstatus_csv_dumper_2667);
    fifo_csv_dumper_2668 = new("./depth2668.csv");
    cstatus_csv_dumper_2668 = new("./chan_status2668.csv");
    fifo_monitor_2668 = new(fifo_csv_dumper_2668,fifo_intf_2668,cstatus_csv_dumper_2668);
    fifo_csv_dumper_2669 = new("./depth2669.csv");
    cstatus_csv_dumper_2669 = new("./chan_status2669.csv");
    fifo_monitor_2669 = new(fifo_csv_dumper_2669,fifo_intf_2669,cstatus_csv_dumper_2669);
    fifo_csv_dumper_2670 = new("./depth2670.csv");
    cstatus_csv_dumper_2670 = new("./chan_status2670.csv");
    fifo_monitor_2670 = new(fifo_csv_dumper_2670,fifo_intf_2670,cstatus_csv_dumper_2670);
    fifo_csv_dumper_2671 = new("./depth2671.csv");
    cstatus_csv_dumper_2671 = new("./chan_status2671.csv");
    fifo_monitor_2671 = new(fifo_csv_dumper_2671,fifo_intf_2671,cstatus_csv_dumper_2671);
    fifo_csv_dumper_2672 = new("./depth2672.csv");
    cstatus_csv_dumper_2672 = new("./chan_status2672.csv");
    fifo_monitor_2672 = new(fifo_csv_dumper_2672,fifo_intf_2672,cstatus_csv_dumper_2672);
    fifo_csv_dumper_2673 = new("./depth2673.csv");
    cstatus_csv_dumper_2673 = new("./chan_status2673.csv");
    fifo_monitor_2673 = new(fifo_csv_dumper_2673,fifo_intf_2673,cstatus_csv_dumper_2673);
    fifo_csv_dumper_2674 = new("./depth2674.csv");
    cstatus_csv_dumper_2674 = new("./chan_status2674.csv");
    fifo_monitor_2674 = new(fifo_csv_dumper_2674,fifo_intf_2674,cstatus_csv_dumper_2674);
    fifo_csv_dumper_2675 = new("./depth2675.csv");
    cstatus_csv_dumper_2675 = new("./chan_status2675.csv");
    fifo_monitor_2675 = new(fifo_csv_dumper_2675,fifo_intf_2675,cstatus_csv_dumper_2675);
    fifo_csv_dumper_2676 = new("./depth2676.csv");
    cstatus_csv_dumper_2676 = new("./chan_status2676.csv");
    fifo_monitor_2676 = new(fifo_csv_dumper_2676,fifo_intf_2676,cstatus_csv_dumper_2676);
    fifo_csv_dumper_2677 = new("./depth2677.csv");
    cstatus_csv_dumper_2677 = new("./chan_status2677.csv");
    fifo_monitor_2677 = new(fifo_csv_dumper_2677,fifo_intf_2677,cstatus_csv_dumper_2677);
    fifo_csv_dumper_2678 = new("./depth2678.csv");
    cstatus_csv_dumper_2678 = new("./chan_status2678.csv");
    fifo_monitor_2678 = new(fifo_csv_dumper_2678,fifo_intf_2678,cstatus_csv_dumper_2678);
    fifo_csv_dumper_2679 = new("./depth2679.csv");
    cstatus_csv_dumper_2679 = new("./chan_status2679.csv");
    fifo_monitor_2679 = new(fifo_csv_dumper_2679,fifo_intf_2679,cstatus_csv_dumper_2679);
    fifo_csv_dumper_2680 = new("./depth2680.csv");
    cstatus_csv_dumper_2680 = new("./chan_status2680.csv");
    fifo_monitor_2680 = new(fifo_csv_dumper_2680,fifo_intf_2680,cstatus_csv_dumper_2680);
    fifo_csv_dumper_2681 = new("./depth2681.csv");
    cstatus_csv_dumper_2681 = new("./chan_status2681.csv");
    fifo_monitor_2681 = new(fifo_csv_dumper_2681,fifo_intf_2681,cstatus_csv_dumper_2681);
    fifo_csv_dumper_2682 = new("./depth2682.csv");
    cstatus_csv_dumper_2682 = new("./chan_status2682.csv");
    fifo_monitor_2682 = new(fifo_csv_dumper_2682,fifo_intf_2682,cstatus_csv_dumper_2682);
    fifo_csv_dumper_2683 = new("./depth2683.csv");
    cstatus_csv_dumper_2683 = new("./chan_status2683.csv");
    fifo_monitor_2683 = new(fifo_csv_dumper_2683,fifo_intf_2683,cstatus_csv_dumper_2683);
    fifo_csv_dumper_2684 = new("./depth2684.csv");
    cstatus_csv_dumper_2684 = new("./chan_status2684.csv");
    fifo_monitor_2684 = new(fifo_csv_dumper_2684,fifo_intf_2684,cstatus_csv_dumper_2684);
    fifo_csv_dumper_2685 = new("./depth2685.csv");
    cstatus_csv_dumper_2685 = new("./chan_status2685.csv");
    fifo_monitor_2685 = new(fifo_csv_dumper_2685,fifo_intf_2685,cstatus_csv_dumper_2685);
    fifo_csv_dumper_2686 = new("./depth2686.csv");
    cstatus_csv_dumper_2686 = new("./chan_status2686.csv");
    fifo_monitor_2686 = new(fifo_csv_dumper_2686,fifo_intf_2686,cstatus_csv_dumper_2686);
    fifo_csv_dumper_2687 = new("./depth2687.csv");
    cstatus_csv_dumper_2687 = new("./chan_status2687.csv");
    fifo_monitor_2687 = new(fifo_csv_dumper_2687,fifo_intf_2687,cstatus_csv_dumper_2687);
    fifo_csv_dumper_2688 = new("./depth2688.csv");
    cstatus_csv_dumper_2688 = new("./chan_status2688.csv");
    fifo_monitor_2688 = new(fifo_csv_dumper_2688,fifo_intf_2688,cstatus_csv_dumper_2688);
    fifo_csv_dumper_2689 = new("./depth2689.csv");
    cstatus_csv_dumper_2689 = new("./chan_status2689.csv");
    fifo_monitor_2689 = new(fifo_csv_dumper_2689,fifo_intf_2689,cstatus_csv_dumper_2689);
    fifo_csv_dumper_2690 = new("./depth2690.csv");
    cstatus_csv_dumper_2690 = new("./chan_status2690.csv");
    fifo_monitor_2690 = new(fifo_csv_dumper_2690,fifo_intf_2690,cstatus_csv_dumper_2690);
    fifo_csv_dumper_2691 = new("./depth2691.csv");
    cstatus_csv_dumper_2691 = new("./chan_status2691.csv");
    fifo_monitor_2691 = new(fifo_csv_dumper_2691,fifo_intf_2691,cstatus_csv_dumper_2691);
    fifo_csv_dumper_2692 = new("./depth2692.csv");
    cstatus_csv_dumper_2692 = new("./chan_status2692.csv");
    fifo_monitor_2692 = new(fifo_csv_dumper_2692,fifo_intf_2692,cstatus_csv_dumper_2692);
    fifo_csv_dumper_2693 = new("./depth2693.csv");
    cstatus_csv_dumper_2693 = new("./chan_status2693.csv");
    fifo_monitor_2693 = new(fifo_csv_dumper_2693,fifo_intf_2693,cstatus_csv_dumper_2693);
    fifo_csv_dumper_2694 = new("./depth2694.csv");
    cstatus_csv_dumper_2694 = new("./chan_status2694.csv");
    fifo_monitor_2694 = new(fifo_csv_dumper_2694,fifo_intf_2694,cstatus_csv_dumper_2694);
    fifo_csv_dumper_2695 = new("./depth2695.csv");
    cstatus_csv_dumper_2695 = new("./chan_status2695.csv");
    fifo_monitor_2695 = new(fifo_csv_dumper_2695,fifo_intf_2695,cstatus_csv_dumper_2695);
    fifo_csv_dumper_2696 = new("./depth2696.csv");
    cstatus_csv_dumper_2696 = new("./chan_status2696.csv");
    fifo_monitor_2696 = new(fifo_csv_dumper_2696,fifo_intf_2696,cstatus_csv_dumper_2696);
    fifo_csv_dumper_2697 = new("./depth2697.csv");
    cstatus_csv_dumper_2697 = new("./chan_status2697.csv");
    fifo_monitor_2697 = new(fifo_csv_dumper_2697,fifo_intf_2697,cstatus_csv_dumper_2697);
    fifo_csv_dumper_2698 = new("./depth2698.csv");
    cstatus_csv_dumper_2698 = new("./chan_status2698.csv");
    fifo_monitor_2698 = new(fifo_csv_dumper_2698,fifo_intf_2698,cstatus_csv_dumper_2698);
    fifo_csv_dumper_2699 = new("./depth2699.csv");
    cstatus_csv_dumper_2699 = new("./chan_status2699.csv");
    fifo_monitor_2699 = new(fifo_csv_dumper_2699,fifo_intf_2699,cstatus_csv_dumper_2699);
    fifo_csv_dumper_2700 = new("./depth2700.csv");
    cstatus_csv_dumper_2700 = new("./chan_status2700.csv");
    fifo_monitor_2700 = new(fifo_csv_dumper_2700,fifo_intf_2700,cstatus_csv_dumper_2700);
    fifo_csv_dumper_2701 = new("./depth2701.csv");
    cstatus_csv_dumper_2701 = new("./chan_status2701.csv");
    fifo_monitor_2701 = new(fifo_csv_dumper_2701,fifo_intf_2701,cstatus_csv_dumper_2701);
    fifo_csv_dumper_2702 = new("./depth2702.csv");
    cstatus_csv_dumper_2702 = new("./chan_status2702.csv");
    fifo_monitor_2702 = new(fifo_csv_dumper_2702,fifo_intf_2702,cstatus_csv_dumper_2702);
    fifo_csv_dumper_2703 = new("./depth2703.csv");
    cstatus_csv_dumper_2703 = new("./chan_status2703.csv");
    fifo_monitor_2703 = new(fifo_csv_dumper_2703,fifo_intf_2703,cstatus_csv_dumper_2703);
    fifo_csv_dumper_2704 = new("./depth2704.csv");
    cstatus_csv_dumper_2704 = new("./chan_status2704.csv");
    fifo_monitor_2704 = new(fifo_csv_dumper_2704,fifo_intf_2704,cstatus_csv_dumper_2704);
    fifo_csv_dumper_2705 = new("./depth2705.csv");
    cstatus_csv_dumper_2705 = new("./chan_status2705.csv");
    fifo_monitor_2705 = new(fifo_csv_dumper_2705,fifo_intf_2705,cstatus_csv_dumper_2705);
    fifo_csv_dumper_2706 = new("./depth2706.csv");
    cstatus_csv_dumper_2706 = new("./chan_status2706.csv");
    fifo_monitor_2706 = new(fifo_csv_dumper_2706,fifo_intf_2706,cstatus_csv_dumper_2706);
    fifo_csv_dumper_2707 = new("./depth2707.csv");
    cstatus_csv_dumper_2707 = new("./chan_status2707.csv");
    fifo_monitor_2707 = new(fifo_csv_dumper_2707,fifo_intf_2707,cstatus_csv_dumper_2707);
    fifo_csv_dumper_2708 = new("./depth2708.csv");
    cstatus_csv_dumper_2708 = new("./chan_status2708.csv");
    fifo_monitor_2708 = new(fifo_csv_dumper_2708,fifo_intf_2708,cstatus_csv_dumper_2708);
    fifo_csv_dumper_2709 = new("./depth2709.csv");
    cstatus_csv_dumper_2709 = new("./chan_status2709.csv");
    fifo_monitor_2709 = new(fifo_csv_dumper_2709,fifo_intf_2709,cstatus_csv_dumper_2709);
    fifo_csv_dumper_2710 = new("./depth2710.csv");
    cstatus_csv_dumper_2710 = new("./chan_status2710.csv");
    fifo_monitor_2710 = new(fifo_csv_dumper_2710,fifo_intf_2710,cstatus_csv_dumper_2710);
    fifo_csv_dumper_2711 = new("./depth2711.csv");
    cstatus_csv_dumper_2711 = new("./chan_status2711.csv");
    fifo_monitor_2711 = new(fifo_csv_dumper_2711,fifo_intf_2711,cstatus_csv_dumper_2711);
    fifo_csv_dumper_2712 = new("./depth2712.csv");
    cstatus_csv_dumper_2712 = new("./chan_status2712.csv");
    fifo_monitor_2712 = new(fifo_csv_dumper_2712,fifo_intf_2712,cstatus_csv_dumper_2712);
    fifo_csv_dumper_2713 = new("./depth2713.csv");
    cstatus_csv_dumper_2713 = new("./chan_status2713.csv");
    fifo_monitor_2713 = new(fifo_csv_dumper_2713,fifo_intf_2713,cstatus_csv_dumper_2713);
    fifo_csv_dumper_2714 = new("./depth2714.csv");
    cstatus_csv_dumper_2714 = new("./chan_status2714.csv");
    fifo_monitor_2714 = new(fifo_csv_dumper_2714,fifo_intf_2714,cstatus_csv_dumper_2714);

    pstall_csv_dumper_1 = new("./stalling1.csv");
    pstatus_csv_dumper_1 = new("./status1.csv");
    process_monitor_1 = new(pstall_csv_dumper_1,process_intf_1,pstatus_csv_dumper_1);
    pstall_csv_dumper_2 = new("./stalling2.csv");
    pstatus_csv_dumper_2 = new("./status2.csv");
    process_monitor_2 = new(pstall_csv_dumper_2,process_intf_2,pstatus_csv_dumper_2);
    pstall_csv_dumper_3 = new("./stalling3.csv");
    pstatus_csv_dumper_3 = new("./status3.csv");
    process_monitor_3 = new(pstall_csv_dumper_3,process_intf_3,pstatus_csv_dumper_3);
    pstall_csv_dumper_4 = new("./stalling4.csv");
    pstatus_csv_dumper_4 = new("./status4.csv");
    process_monitor_4 = new(pstall_csv_dumper_4,process_intf_4,pstatus_csv_dumper_4);

    mstatus_csv_dumper_1 = new("./module_status1.csv");
    module_monitor_1 = new(module_intf_1,mstatus_csv_dumper_1);
    mstatus_csv_dumper_2 = new("./module_status2.csv");
    module_monitor_2 = new(module_intf_2,mstatus_csv_dumper_2);
    mstatus_csv_dumper_3 = new("./module_status3.csv");
    module_monitor_3 = new(module_intf_3,mstatus_csv_dumper_3);



    seq_loop_csv_dumper_1 = new("./seq_loop_status1.csv");
    seq_loop_monitor_1 = new(seq_loop_intf_1,seq_loop_csv_dumper_1);

    upc_loop_csv_dumper_1 = new("./upc_loop_status1.csv");
    upc_loop_monitor_1 = new(upc_loop_intf_1,upc_loop_csv_dumper_1);

    sample_manager_inst.add_one_monitor(fifo_monitor_1);
    sample_manager_inst.add_one_monitor(fifo_monitor_2);
    sample_manager_inst.add_one_monitor(fifo_monitor_3);
    sample_manager_inst.add_one_monitor(fifo_monitor_4);
    sample_manager_inst.add_one_monitor(fifo_monitor_5);
    sample_manager_inst.add_one_monitor(fifo_monitor_6);
    sample_manager_inst.add_one_monitor(fifo_monitor_7);
    sample_manager_inst.add_one_monitor(fifo_monitor_8);
    sample_manager_inst.add_one_monitor(fifo_monitor_9);
    sample_manager_inst.add_one_monitor(fifo_monitor_10);
    sample_manager_inst.add_one_monitor(fifo_monitor_11);
    sample_manager_inst.add_one_monitor(fifo_monitor_12);
    sample_manager_inst.add_one_monitor(fifo_monitor_13);
    sample_manager_inst.add_one_monitor(fifo_monitor_14);
    sample_manager_inst.add_one_monitor(fifo_monitor_15);
    sample_manager_inst.add_one_monitor(fifo_monitor_16);
    sample_manager_inst.add_one_monitor(fifo_monitor_17);
    sample_manager_inst.add_one_monitor(fifo_monitor_18);
    sample_manager_inst.add_one_monitor(fifo_monitor_19);
    sample_manager_inst.add_one_monitor(fifo_monitor_20);
    sample_manager_inst.add_one_monitor(fifo_monitor_21);
    sample_manager_inst.add_one_monitor(fifo_monitor_22);
    sample_manager_inst.add_one_monitor(fifo_monitor_23);
    sample_manager_inst.add_one_monitor(fifo_monitor_24);
    sample_manager_inst.add_one_monitor(fifo_monitor_25);
    sample_manager_inst.add_one_monitor(fifo_monitor_26);
    sample_manager_inst.add_one_monitor(fifo_monitor_27);
    sample_manager_inst.add_one_monitor(fifo_monitor_28);
    sample_manager_inst.add_one_monitor(fifo_monitor_29);
    sample_manager_inst.add_one_monitor(fifo_monitor_30);
    sample_manager_inst.add_one_monitor(fifo_monitor_31);
    sample_manager_inst.add_one_monitor(fifo_monitor_32);
    sample_manager_inst.add_one_monitor(fifo_monitor_33);
    sample_manager_inst.add_one_monitor(fifo_monitor_34);
    sample_manager_inst.add_one_monitor(fifo_monitor_35);
    sample_manager_inst.add_one_monitor(fifo_monitor_36);
    sample_manager_inst.add_one_monitor(fifo_monitor_37);
    sample_manager_inst.add_one_monitor(fifo_monitor_38);
    sample_manager_inst.add_one_monitor(fifo_monitor_39);
    sample_manager_inst.add_one_monitor(fifo_monitor_40);
    sample_manager_inst.add_one_monitor(fifo_monitor_41);
    sample_manager_inst.add_one_monitor(fifo_monitor_42);
    sample_manager_inst.add_one_monitor(fifo_monitor_43);
    sample_manager_inst.add_one_monitor(fifo_monitor_44);
    sample_manager_inst.add_one_monitor(fifo_monitor_45);
    sample_manager_inst.add_one_monitor(fifo_monitor_46);
    sample_manager_inst.add_one_monitor(fifo_monitor_47);
    sample_manager_inst.add_one_monitor(fifo_monitor_48);
    sample_manager_inst.add_one_monitor(fifo_monitor_49);
    sample_manager_inst.add_one_monitor(fifo_monitor_50);
    sample_manager_inst.add_one_monitor(fifo_monitor_51);
    sample_manager_inst.add_one_monitor(fifo_monitor_52);
    sample_manager_inst.add_one_monitor(fifo_monitor_53);
    sample_manager_inst.add_one_monitor(fifo_monitor_54);
    sample_manager_inst.add_one_monitor(fifo_monitor_55);
    sample_manager_inst.add_one_monitor(fifo_monitor_56);
    sample_manager_inst.add_one_monitor(fifo_monitor_57);
    sample_manager_inst.add_one_monitor(fifo_monitor_58);
    sample_manager_inst.add_one_monitor(fifo_monitor_59);
    sample_manager_inst.add_one_monitor(fifo_monitor_60);
    sample_manager_inst.add_one_monitor(fifo_monitor_61);
    sample_manager_inst.add_one_monitor(fifo_monitor_62);
    sample_manager_inst.add_one_monitor(fifo_monitor_63);
    sample_manager_inst.add_one_monitor(fifo_monitor_64);
    sample_manager_inst.add_one_monitor(fifo_monitor_65);
    sample_manager_inst.add_one_monitor(fifo_monitor_66);
    sample_manager_inst.add_one_monitor(fifo_monitor_67);
    sample_manager_inst.add_one_monitor(fifo_monitor_68);
    sample_manager_inst.add_one_monitor(fifo_monitor_69);
    sample_manager_inst.add_one_monitor(fifo_monitor_70);
    sample_manager_inst.add_one_monitor(fifo_monitor_71);
    sample_manager_inst.add_one_monitor(fifo_monitor_72);
    sample_manager_inst.add_one_monitor(fifo_monitor_73);
    sample_manager_inst.add_one_monitor(fifo_monitor_74);
    sample_manager_inst.add_one_monitor(fifo_monitor_75);
    sample_manager_inst.add_one_monitor(fifo_monitor_76);
    sample_manager_inst.add_one_monitor(fifo_monitor_77);
    sample_manager_inst.add_one_monitor(fifo_monitor_78);
    sample_manager_inst.add_one_monitor(fifo_monitor_79);
    sample_manager_inst.add_one_monitor(fifo_monitor_80);
    sample_manager_inst.add_one_monitor(fifo_monitor_81);
    sample_manager_inst.add_one_monitor(fifo_monitor_82);
    sample_manager_inst.add_one_monitor(fifo_monitor_83);
    sample_manager_inst.add_one_monitor(fifo_monitor_84);
    sample_manager_inst.add_one_monitor(fifo_monitor_85);
    sample_manager_inst.add_one_monitor(fifo_monitor_86);
    sample_manager_inst.add_one_monitor(fifo_monitor_87);
    sample_manager_inst.add_one_monitor(fifo_monitor_88);
    sample_manager_inst.add_one_monitor(fifo_monitor_89);
    sample_manager_inst.add_one_monitor(fifo_monitor_90);
    sample_manager_inst.add_one_monitor(fifo_monitor_91);
    sample_manager_inst.add_one_monitor(fifo_monitor_92);
    sample_manager_inst.add_one_monitor(fifo_monitor_93);
    sample_manager_inst.add_one_monitor(fifo_monitor_94);
    sample_manager_inst.add_one_monitor(fifo_monitor_95);
    sample_manager_inst.add_one_monitor(fifo_monitor_96);
    sample_manager_inst.add_one_monitor(fifo_monitor_97);
    sample_manager_inst.add_one_monitor(fifo_monitor_98);
    sample_manager_inst.add_one_monitor(fifo_monitor_99);
    sample_manager_inst.add_one_monitor(fifo_monitor_100);
    sample_manager_inst.add_one_monitor(fifo_monitor_101);
    sample_manager_inst.add_one_monitor(fifo_monitor_102);
    sample_manager_inst.add_one_monitor(fifo_monitor_103);
    sample_manager_inst.add_one_monitor(fifo_monitor_104);
    sample_manager_inst.add_one_monitor(fifo_monitor_105);
    sample_manager_inst.add_one_monitor(fifo_monitor_106);
    sample_manager_inst.add_one_monitor(fifo_monitor_107);
    sample_manager_inst.add_one_monitor(fifo_monitor_108);
    sample_manager_inst.add_one_monitor(fifo_monitor_109);
    sample_manager_inst.add_one_monitor(fifo_monitor_110);
    sample_manager_inst.add_one_monitor(fifo_monitor_111);
    sample_manager_inst.add_one_monitor(fifo_monitor_112);
    sample_manager_inst.add_one_monitor(fifo_monitor_113);
    sample_manager_inst.add_one_monitor(fifo_monitor_114);
    sample_manager_inst.add_one_monitor(fifo_monitor_115);
    sample_manager_inst.add_one_monitor(fifo_monitor_116);
    sample_manager_inst.add_one_monitor(fifo_monitor_117);
    sample_manager_inst.add_one_monitor(fifo_monitor_118);
    sample_manager_inst.add_one_monitor(fifo_monitor_119);
    sample_manager_inst.add_one_monitor(fifo_monitor_120);
    sample_manager_inst.add_one_monitor(fifo_monitor_121);
    sample_manager_inst.add_one_monitor(fifo_monitor_122);
    sample_manager_inst.add_one_monitor(fifo_monitor_123);
    sample_manager_inst.add_one_monitor(fifo_monitor_124);
    sample_manager_inst.add_one_monitor(fifo_monitor_125);
    sample_manager_inst.add_one_monitor(fifo_monitor_126);
    sample_manager_inst.add_one_monitor(fifo_monitor_127);
    sample_manager_inst.add_one_monitor(fifo_monitor_128);
    sample_manager_inst.add_one_monitor(fifo_monitor_129);
    sample_manager_inst.add_one_monitor(fifo_monitor_130);
    sample_manager_inst.add_one_monitor(fifo_monitor_131);
    sample_manager_inst.add_one_monitor(fifo_monitor_132);
    sample_manager_inst.add_one_monitor(fifo_monitor_133);
    sample_manager_inst.add_one_monitor(fifo_monitor_134);
    sample_manager_inst.add_one_monitor(fifo_monitor_135);
    sample_manager_inst.add_one_monitor(fifo_monitor_136);
    sample_manager_inst.add_one_monitor(fifo_monitor_137);
    sample_manager_inst.add_one_monitor(fifo_monitor_138);
    sample_manager_inst.add_one_monitor(fifo_monitor_139);
    sample_manager_inst.add_one_monitor(fifo_monitor_140);
    sample_manager_inst.add_one_monitor(fifo_monitor_141);
    sample_manager_inst.add_one_monitor(fifo_monitor_142);
    sample_manager_inst.add_one_monitor(fifo_monitor_143);
    sample_manager_inst.add_one_monitor(fifo_monitor_144);
    sample_manager_inst.add_one_monitor(fifo_monitor_145);
    sample_manager_inst.add_one_monitor(fifo_monitor_146);
    sample_manager_inst.add_one_monitor(fifo_monitor_147);
    sample_manager_inst.add_one_monitor(fifo_monitor_148);
    sample_manager_inst.add_one_monitor(fifo_monitor_149);
    sample_manager_inst.add_one_monitor(fifo_monitor_150);
    sample_manager_inst.add_one_monitor(fifo_monitor_151);
    sample_manager_inst.add_one_monitor(fifo_monitor_152);
    sample_manager_inst.add_one_monitor(fifo_monitor_153);
    sample_manager_inst.add_one_monitor(fifo_monitor_154);
    sample_manager_inst.add_one_monitor(fifo_monitor_155);
    sample_manager_inst.add_one_monitor(fifo_monitor_156);
    sample_manager_inst.add_one_monitor(fifo_monitor_157);
    sample_manager_inst.add_one_monitor(fifo_monitor_158);
    sample_manager_inst.add_one_monitor(fifo_monitor_159);
    sample_manager_inst.add_one_monitor(fifo_monitor_160);
    sample_manager_inst.add_one_monitor(fifo_monitor_161);
    sample_manager_inst.add_one_monitor(fifo_monitor_162);
    sample_manager_inst.add_one_monitor(fifo_monitor_163);
    sample_manager_inst.add_one_monitor(fifo_monitor_164);
    sample_manager_inst.add_one_monitor(fifo_monitor_165);
    sample_manager_inst.add_one_monitor(fifo_monitor_166);
    sample_manager_inst.add_one_monitor(fifo_monitor_167);
    sample_manager_inst.add_one_monitor(fifo_monitor_168);
    sample_manager_inst.add_one_monitor(fifo_monitor_169);
    sample_manager_inst.add_one_monitor(fifo_monitor_170);
    sample_manager_inst.add_one_monitor(fifo_monitor_171);
    sample_manager_inst.add_one_monitor(fifo_monitor_172);
    sample_manager_inst.add_one_monitor(fifo_monitor_173);
    sample_manager_inst.add_one_monitor(fifo_monitor_174);
    sample_manager_inst.add_one_monitor(fifo_monitor_175);
    sample_manager_inst.add_one_monitor(fifo_monitor_176);
    sample_manager_inst.add_one_monitor(fifo_monitor_177);
    sample_manager_inst.add_one_monitor(fifo_monitor_178);
    sample_manager_inst.add_one_monitor(fifo_monitor_179);
    sample_manager_inst.add_one_monitor(fifo_monitor_180);
    sample_manager_inst.add_one_monitor(fifo_monitor_181);
    sample_manager_inst.add_one_monitor(fifo_monitor_182);
    sample_manager_inst.add_one_monitor(fifo_monitor_183);
    sample_manager_inst.add_one_monitor(fifo_monitor_184);
    sample_manager_inst.add_one_monitor(fifo_monitor_185);
    sample_manager_inst.add_one_monitor(fifo_monitor_186);
    sample_manager_inst.add_one_monitor(fifo_monitor_187);
    sample_manager_inst.add_one_monitor(fifo_monitor_188);
    sample_manager_inst.add_one_monitor(fifo_monitor_189);
    sample_manager_inst.add_one_monitor(fifo_monitor_190);
    sample_manager_inst.add_one_monitor(fifo_monitor_191);
    sample_manager_inst.add_one_monitor(fifo_monitor_192);
    sample_manager_inst.add_one_monitor(fifo_monitor_193);
    sample_manager_inst.add_one_monitor(fifo_monitor_194);
    sample_manager_inst.add_one_monitor(fifo_monitor_195);
    sample_manager_inst.add_one_monitor(fifo_monitor_196);
    sample_manager_inst.add_one_monitor(fifo_monitor_197);
    sample_manager_inst.add_one_monitor(fifo_monitor_198);
    sample_manager_inst.add_one_monitor(fifo_monitor_199);
    sample_manager_inst.add_one_monitor(fifo_monitor_200);
    sample_manager_inst.add_one_monitor(fifo_monitor_201);
    sample_manager_inst.add_one_monitor(fifo_monitor_202);
    sample_manager_inst.add_one_monitor(fifo_monitor_203);
    sample_manager_inst.add_one_monitor(fifo_monitor_204);
    sample_manager_inst.add_one_monitor(fifo_monitor_205);
    sample_manager_inst.add_one_monitor(fifo_monitor_206);
    sample_manager_inst.add_one_monitor(fifo_monitor_207);
    sample_manager_inst.add_one_monitor(fifo_monitor_208);
    sample_manager_inst.add_one_monitor(fifo_monitor_209);
    sample_manager_inst.add_one_monitor(fifo_monitor_210);
    sample_manager_inst.add_one_monitor(fifo_monitor_211);
    sample_manager_inst.add_one_monitor(fifo_monitor_212);
    sample_manager_inst.add_one_monitor(fifo_monitor_213);
    sample_manager_inst.add_one_monitor(fifo_monitor_214);
    sample_manager_inst.add_one_monitor(fifo_monitor_215);
    sample_manager_inst.add_one_monitor(fifo_monitor_216);
    sample_manager_inst.add_one_monitor(fifo_monitor_217);
    sample_manager_inst.add_one_monitor(fifo_monitor_218);
    sample_manager_inst.add_one_monitor(fifo_monitor_219);
    sample_manager_inst.add_one_monitor(fifo_monitor_220);
    sample_manager_inst.add_one_monitor(fifo_monitor_221);
    sample_manager_inst.add_one_monitor(fifo_monitor_222);
    sample_manager_inst.add_one_monitor(fifo_monitor_223);
    sample_manager_inst.add_one_monitor(fifo_monitor_224);
    sample_manager_inst.add_one_monitor(fifo_monitor_225);
    sample_manager_inst.add_one_monitor(fifo_monitor_226);
    sample_manager_inst.add_one_monitor(fifo_monitor_227);
    sample_manager_inst.add_one_monitor(fifo_monitor_228);
    sample_manager_inst.add_one_monitor(fifo_monitor_229);
    sample_manager_inst.add_one_monitor(fifo_monitor_230);
    sample_manager_inst.add_one_monitor(fifo_monitor_231);
    sample_manager_inst.add_one_monitor(fifo_monitor_232);
    sample_manager_inst.add_one_monitor(fifo_monitor_233);
    sample_manager_inst.add_one_monitor(fifo_monitor_234);
    sample_manager_inst.add_one_monitor(fifo_monitor_235);
    sample_manager_inst.add_one_monitor(fifo_monitor_236);
    sample_manager_inst.add_one_monitor(fifo_monitor_237);
    sample_manager_inst.add_one_monitor(fifo_monitor_238);
    sample_manager_inst.add_one_monitor(fifo_monitor_239);
    sample_manager_inst.add_one_monitor(fifo_monitor_240);
    sample_manager_inst.add_one_monitor(fifo_monitor_241);
    sample_manager_inst.add_one_monitor(fifo_monitor_242);
    sample_manager_inst.add_one_monitor(fifo_monitor_243);
    sample_manager_inst.add_one_monitor(fifo_monitor_244);
    sample_manager_inst.add_one_monitor(fifo_monitor_245);
    sample_manager_inst.add_one_monitor(fifo_monitor_246);
    sample_manager_inst.add_one_monitor(fifo_monitor_247);
    sample_manager_inst.add_one_monitor(fifo_monitor_248);
    sample_manager_inst.add_one_monitor(fifo_monitor_249);
    sample_manager_inst.add_one_monitor(fifo_monitor_250);
    sample_manager_inst.add_one_monitor(fifo_monitor_251);
    sample_manager_inst.add_one_monitor(fifo_monitor_252);
    sample_manager_inst.add_one_monitor(fifo_monitor_253);
    sample_manager_inst.add_one_monitor(fifo_monitor_254);
    sample_manager_inst.add_one_monitor(fifo_monitor_255);
    sample_manager_inst.add_one_monitor(fifo_monitor_256);
    sample_manager_inst.add_one_monitor(fifo_monitor_257);
    sample_manager_inst.add_one_monitor(fifo_monitor_258);
    sample_manager_inst.add_one_monitor(fifo_monitor_259);
    sample_manager_inst.add_one_monitor(fifo_monitor_260);
    sample_manager_inst.add_one_monitor(fifo_monitor_261);
    sample_manager_inst.add_one_monitor(fifo_monitor_262);
    sample_manager_inst.add_one_monitor(fifo_monitor_263);
    sample_manager_inst.add_one_monitor(fifo_monitor_264);
    sample_manager_inst.add_one_monitor(fifo_monitor_265);
    sample_manager_inst.add_one_monitor(fifo_monitor_266);
    sample_manager_inst.add_one_monitor(fifo_monitor_267);
    sample_manager_inst.add_one_monitor(fifo_monitor_268);
    sample_manager_inst.add_one_monitor(fifo_monitor_269);
    sample_manager_inst.add_one_monitor(fifo_monitor_270);
    sample_manager_inst.add_one_monitor(fifo_monitor_271);
    sample_manager_inst.add_one_monitor(fifo_monitor_272);
    sample_manager_inst.add_one_monitor(fifo_monitor_273);
    sample_manager_inst.add_one_monitor(fifo_monitor_274);
    sample_manager_inst.add_one_monitor(fifo_monitor_275);
    sample_manager_inst.add_one_monitor(fifo_monitor_276);
    sample_manager_inst.add_one_monitor(fifo_monitor_277);
    sample_manager_inst.add_one_monitor(fifo_monitor_278);
    sample_manager_inst.add_one_monitor(fifo_monitor_279);
    sample_manager_inst.add_one_monitor(fifo_monitor_280);
    sample_manager_inst.add_one_monitor(fifo_monitor_281);
    sample_manager_inst.add_one_monitor(fifo_monitor_282);
    sample_manager_inst.add_one_monitor(fifo_monitor_283);
    sample_manager_inst.add_one_monitor(fifo_monitor_284);
    sample_manager_inst.add_one_monitor(fifo_monitor_285);
    sample_manager_inst.add_one_monitor(fifo_monitor_286);
    sample_manager_inst.add_one_monitor(fifo_monitor_287);
    sample_manager_inst.add_one_monitor(fifo_monitor_288);
    sample_manager_inst.add_one_monitor(fifo_monitor_289);
    sample_manager_inst.add_one_monitor(fifo_monitor_290);
    sample_manager_inst.add_one_monitor(fifo_monitor_291);
    sample_manager_inst.add_one_monitor(fifo_monitor_292);
    sample_manager_inst.add_one_monitor(fifo_monitor_293);
    sample_manager_inst.add_one_monitor(fifo_monitor_294);
    sample_manager_inst.add_one_monitor(fifo_monitor_295);
    sample_manager_inst.add_one_monitor(fifo_monitor_296);
    sample_manager_inst.add_one_monitor(fifo_monitor_297);
    sample_manager_inst.add_one_monitor(fifo_monitor_298);
    sample_manager_inst.add_one_monitor(fifo_monitor_299);
    sample_manager_inst.add_one_monitor(fifo_monitor_300);
    sample_manager_inst.add_one_monitor(fifo_monitor_301);
    sample_manager_inst.add_one_monitor(fifo_monitor_302);
    sample_manager_inst.add_one_monitor(fifo_monitor_303);
    sample_manager_inst.add_one_monitor(fifo_monitor_304);
    sample_manager_inst.add_one_monitor(fifo_monitor_305);
    sample_manager_inst.add_one_monitor(fifo_monitor_306);
    sample_manager_inst.add_one_monitor(fifo_monitor_307);
    sample_manager_inst.add_one_monitor(fifo_monitor_308);
    sample_manager_inst.add_one_monitor(fifo_monitor_309);
    sample_manager_inst.add_one_monitor(fifo_monitor_310);
    sample_manager_inst.add_one_monitor(fifo_monitor_311);
    sample_manager_inst.add_one_monitor(fifo_monitor_312);
    sample_manager_inst.add_one_monitor(fifo_monitor_313);
    sample_manager_inst.add_one_monitor(fifo_monitor_314);
    sample_manager_inst.add_one_monitor(fifo_monitor_315);
    sample_manager_inst.add_one_monitor(fifo_monitor_316);
    sample_manager_inst.add_one_monitor(fifo_monitor_317);
    sample_manager_inst.add_one_monitor(fifo_monitor_318);
    sample_manager_inst.add_one_monitor(fifo_monitor_319);
    sample_manager_inst.add_one_monitor(fifo_monitor_320);
    sample_manager_inst.add_one_monitor(fifo_monitor_321);
    sample_manager_inst.add_one_monitor(fifo_monitor_322);
    sample_manager_inst.add_one_monitor(fifo_monitor_323);
    sample_manager_inst.add_one_monitor(fifo_monitor_324);
    sample_manager_inst.add_one_monitor(fifo_monitor_325);
    sample_manager_inst.add_one_monitor(fifo_monitor_326);
    sample_manager_inst.add_one_monitor(fifo_monitor_327);
    sample_manager_inst.add_one_monitor(fifo_monitor_328);
    sample_manager_inst.add_one_monitor(fifo_monitor_329);
    sample_manager_inst.add_one_monitor(fifo_monitor_330);
    sample_manager_inst.add_one_monitor(fifo_monitor_331);
    sample_manager_inst.add_one_monitor(fifo_monitor_332);
    sample_manager_inst.add_one_monitor(fifo_monitor_333);
    sample_manager_inst.add_one_monitor(fifo_monitor_334);
    sample_manager_inst.add_one_monitor(fifo_monitor_335);
    sample_manager_inst.add_one_monitor(fifo_monitor_336);
    sample_manager_inst.add_one_monitor(fifo_monitor_337);
    sample_manager_inst.add_one_monitor(fifo_monitor_338);
    sample_manager_inst.add_one_monitor(fifo_monitor_339);
    sample_manager_inst.add_one_monitor(fifo_monitor_340);
    sample_manager_inst.add_one_monitor(fifo_monitor_341);
    sample_manager_inst.add_one_monitor(fifo_monitor_342);
    sample_manager_inst.add_one_monitor(fifo_monitor_343);
    sample_manager_inst.add_one_monitor(fifo_monitor_344);
    sample_manager_inst.add_one_monitor(fifo_monitor_345);
    sample_manager_inst.add_one_monitor(fifo_monitor_346);
    sample_manager_inst.add_one_monitor(fifo_monitor_347);
    sample_manager_inst.add_one_monitor(fifo_monitor_348);
    sample_manager_inst.add_one_monitor(fifo_monitor_349);
    sample_manager_inst.add_one_monitor(fifo_monitor_350);
    sample_manager_inst.add_one_monitor(fifo_monitor_351);
    sample_manager_inst.add_one_monitor(fifo_monitor_352);
    sample_manager_inst.add_one_monitor(fifo_monitor_353);
    sample_manager_inst.add_one_monitor(fifo_monitor_354);
    sample_manager_inst.add_one_monitor(fifo_monitor_355);
    sample_manager_inst.add_one_monitor(fifo_monitor_356);
    sample_manager_inst.add_one_monitor(fifo_monitor_357);
    sample_manager_inst.add_one_monitor(fifo_monitor_358);
    sample_manager_inst.add_one_monitor(fifo_monitor_359);
    sample_manager_inst.add_one_monitor(fifo_monitor_360);
    sample_manager_inst.add_one_monitor(fifo_monitor_361);
    sample_manager_inst.add_one_monitor(fifo_monitor_362);
    sample_manager_inst.add_one_monitor(fifo_monitor_363);
    sample_manager_inst.add_one_monitor(fifo_monitor_364);
    sample_manager_inst.add_one_monitor(fifo_monitor_365);
    sample_manager_inst.add_one_monitor(fifo_monitor_366);
    sample_manager_inst.add_one_monitor(fifo_monitor_367);
    sample_manager_inst.add_one_monitor(fifo_monitor_368);
    sample_manager_inst.add_one_monitor(fifo_monitor_369);
    sample_manager_inst.add_one_monitor(fifo_monitor_370);
    sample_manager_inst.add_one_monitor(fifo_monitor_371);
    sample_manager_inst.add_one_monitor(fifo_monitor_372);
    sample_manager_inst.add_one_monitor(fifo_monitor_373);
    sample_manager_inst.add_one_monitor(fifo_monitor_374);
    sample_manager_inst.add_one_monitor(fifo_monitor_375);
    sample_manager_inst.add_one_monitor(fifo_monitor_376);
    sample_manager_inst.add_one_monitor(fifo_monitor_377);
    sample_manager_inst.add_one_monitor(fifo_monitor_378);
    sample_manager_inst.add_one_monitor(fifo_monitor_379);
    sample_manager_inst.add_one_monitor(fifo_monitor_380);
    sample_manager_inst.add_one_monitor(fifo_monitor_381);
    sample_manager_inst.add_one_monitor(fifo_monitor_382);
    sample_manager_inst.add_one_monitor(fifo_monitor_383);
    sample_manager_inst.add_one_monitor(fifo_monitor_384);
    sample_manager_inst.add_one_monitor(fifo_monitor_385);
    sample_manager_inst.add_one_monitor(fifo_monitor_386);
    sample_manager_inst.add_one_monitor(fifo_monitor_387);
    sample_manager_inst.add_one_monitor(fifo_monitor_388);
    sample_manager_inst.add_one_monitor(fifo_monitor_389);
    sample_manager_inst.add_one_monitor(fifo_monitor_390);
    sample_manager_inst.add_one_monitor(fifo_monitor_391);
    sample_manager_inst.add_one_monitor(fifo_monitor_392);
    sample_manager_inst.add_one_monitor(fifo_monitor_393);
    sample_manager_inst.add_one_monitor(fifo_monitor_394);
    sample_manager_inst.add_one_monitor(fifo_monitor_395);
    sample_manager_inst.add_one_monitor(fifo_monitor_396);
    sample_manager_inst.add_one_monitor(fifo_monitor_397);
    sample_manager_inst.add_one_monitor(fifo_monitor_398);
    sample_manager_inst.add_one_monitor(fifo_monitor_399);
    sample_manager_inst.add_one_monitor(fifo_monitor_400);
    sample_manager_inst.add_one_monitor(fifo_monitor_401);
    sample_manager_inst.add_one_monitor(fifo_monitor_402);
    sample_manager_inst.add_one_monitor(fifo_monitor_403);
    sample_manager_inst.add_one_monitor(fifo_monitor_404);
    sample_manager_inst.add_one_monitor(fifo_monitor_405);
    sample_manager_inst.add_one_monitor(fifo_monitor_406);
    sample_manager_inst.add_one_monitor(fifo_monitor_407);
    sample_manager_inst.add_one_monitor(fifo_monitor_408);
    sample_manager_inst.add_one_monitor(fifo_monitor_409);
    sample_manager_inst.add_one_monitor(fifo_monitor_410);
    sample_manager_inst.add_one_monitor(fifo_monitor_411);
    sample_manager_inst.add_one_monitor(fifo_monitor_412);
    sample_manager_inst.add_one_monitor(fifo_monitor_413);
    sample_manager_inst.add_one_monitor(fifo_monitor_414);
    sample_manager_inst.add_one_monitor(fifo_monitor_415);
    sample_manager_inst.add_one_monitor(fifo_monitor_416);
    sample_manager_inst.add_one_monitor(fifo_monitor_417);
    sample_manager_inst.add_one_monitor(fifo_monitor_418);
    sample_manager_inst.add_one_monitor(fifo_monitor_419);
    sample_manager_inst.add_one_monitor(fifo_monitor_420);
    sample_manager_inst.add_one_monitor(fifo_monitor_421);
    sample_manager_inst.add_one_monitor(fifo_monitor_422);
    sample_manager_inst.add_one_monitor(fifo_monitor_423);
    sample_manager_inst.add_one_monitor(fifo_monitor_424);
    sample_manager_inst.add_one_monitor(fifo_monitor_425);
    sample_manager_inst.add_one_monitor(fifo_monitor_426);
    sample_manager_inst.add_one_monitor(fifo_monitor_427);
    sample_manager_inst.add_one_monitor(fifo_monitor_428);
    sample_manager_inst.add_one_monitor(fifo_monitor_429);
    sample_manager_inst.add_one_monitor(fifo_monitor_430);
    sample_manager_inst.add_one_monitor(fifo_monitor_431);
    sample_manager_inst.add_one_monitor(fifo_monitor_432);
    sample_manager_inst.add_one_monitor(fifo_monitor_433);
    sample_manager_inst.add_one_monitor(fifo_monitor_434);
    sample_manager_inst.add_one_monitor(fifo_monitor_435);
    sample_manager_inst.add_one_monitor(fifo_monitor_436);
    sample_manager_inst.add_one_monitor(fifo_monitor_437);
    sample_manager_inst.add_one_monitor(fifo_monitor_438);
    sample_manager_inst.add_one_monitor(fifo_monitor_439);
    sample_manager_inst.add_one_monitor(fifo_monitor_440);
    sample_manager_inst.add_one_monitor(fifo_monitor_441);
    sample_manager_inst.add_one_monitor(fifo_monitor_442);
    sample_manager_inst.add_one_monitor(fifo_monitor_443);
    sample_manager_inst.add_one_monitor(fifo_monitor_444);
    sample_manager_inst.add_one_monitor(fifo_monitor_445);
    sample_manager_inst.add_one_monitor(fifo_monitor_446);
    sample_manager_inst.add_one_monitor(fifo_monitor_447);
    sample_manager_inst.add_one_monitor(fifo_monitor_448);
    sample_manager_inst.add_one_monitor(fifo_monitor_449);
    sample_manager_inst.add_one_monitor(fifo_monitor_450);
    sample_manager_inst.add_one_monitor(fifo_monitor_451);
    sample_manager_inst.add_one_monitor(fifo_monitor_452);
    sample_manager_inst.add_one_monitor(fifo_monitor_453);
    sample_manager_inst.add_one_monitor(fifo_monitor_454);
    sample_manager_inst.add_one_monitor(fifo_monitor_455);
    sample_manager_inst.add_one_monitor(fifo_monitor_456);
    sample_manager_inst.add_one_monitor(fifo_monitor_457);
    sample_manager_inst.add_one_monitor(fifo_monitor_458);
    sample_manager_inst.add_one_monitor(fifo_monitor_459);
    sample_manager_inst.add_one_monitor(fifo_monitor_460);
    sample_manager_inst.add_one_monitor(fifo_monitor_461);
    sample_manager_inst.add_one_monitor(fifo_monitor_462);
    sample_manager_inst.add_one_monitor(fifo_monitor_463);
    sample_manager_inst.add_one_monitor(fifo_monitor_464);
    sample_manager_inst.add_one_monitor(fifo_monitor_465);
    sample_manager_inst.add_one_monitor(fifo_monitor_466);
    sample_manager_inst.add_one_monitor(fifo_monitor_467);
    sample_manager_inst.add_one_monitor(fifo_monitor_468);
    sample_manager_inst.add_one_monitor(fifo_monitor_469);
    sample_manager_inst.add_one_monitor(fifo_monitor_470);
    sample_manager_inst.add_one_monitor(fifo_monitor_471);
    sample_manager_inst.add_one_monitor(fifo_monitor_472);
    sample_manager_inst.add_one_monitor(fifo_monitor_473);
    sample_manager_inst.add_one_monitor(fifo_monitor_474);
    sample_manager_inst.add_one_monitor(fifo_monitor_475);
    sample_manager_inst.add_one_monitor(fifo_monitor_476);
    sample_manager_inst.add_one_monitor(fifo_monitor_477);
    sample_manager_inst.add_one_monitor(fifo_monitor_478);
    sample_manager_inst.add_one_monitor(fifo_monitor_479);
    sample_manager_inst.add_one_monitor(fifo_monitor_480);
    sample_manager_inst.add_one_monitor(fifo_monitor_481);
    sample_manager_inst.add_one_monitor(fifo_monitor_482);
    sample_manager_inst.add_one_monitor(fifo_monitor_483);
    sample_manager_inst.add_one_monitor(fifo_monitor_484);
    sample_manager_inst.add_one_monitor(fifo_monitor_485);
    sample_manager_inst.add_one_monitor(fifo_monitor_486);
    sample_manager_inst.add_one_monitor(fifo_monitor_487);
    sample_manager_inst.add_one_monitor(fifo_monitor_488);
    sample_manager_inst.add_one_monitor(fifo_monitor_489);
    sample_manager_inst.add_one_monitor(fifo_monitor_490);
    sample_manager_inst.add_one_monitor(fifo_monitor_491);
    sample_manager_inst.add_one_monitor(fifo_monitor_492);
    sample_manager_inst.add_one_monitor(fifo_monitor_493);
    sample_manager_inst.add_one_monitor(fifo_monitor_494);
    sample_manager_inst.add_one_monitor(fifo_monitor_495);
    sample_manager_inst.add_one_monitor(fifo_monitor_496);
    sample_manager_inst.add_one_monitor(fifo_monitor_497);
    sample_manager_inst.add_one_monitor(fifo_monitor_498);
    sample_manager_inst.add_one_monitor(fifo_monitor_499);
    sample_manager_inst.add_one_monitor(fifo_monitor_500);
    sample_manager_inst.add_one_monitor(fifo_monitor_501);
    sample_manager_inst.add_one_monitor(fifo_monitor_502);
    sample_manager_inst.add_one_monitor(fifo_monitor_503);
    sample_manager_inst.add_one_monitor(fifo_monitor_504);
    sample_manager_inst.add_one_monitor(fifo_monitor_505);
    sample_manager_inst.add_one_monitor(fifo_monitor_506);
    sample_manager_inst.add_one_monitor(fifo_monitor_507);
    sample_manager_inst.add_one_monitor(fifo_monitor_508);
    sample_manager_inst.add_one_monitor(fifo_monitor_509);
    sample_manager_inst.add_one_monitor(fifo_monitor_510);
    sample_manager_inst.add_one_monitor(fifo_monitor_511);
    sample_manager_inst.add_one_monitor(fifo_monitor_512);
    sample_manager_inst.add_one_monitor(fifo_monitor_513);
    sample_manager_inst.add_one_monitor(fifo_monitor_514);
    sample_manager_inst.add_one_monitor(fifo_monitor_515);
    sample_manager_inst.add_one_monitor(fifo_monitor_516);
    sample_manager_inst.add_one_monitor(fifo_monitor_517);
    sample_manager_inst.add_one_monitor(fifo_monitor_518);
    sample_manager_inst.add_one_monitor(fifo_monitor_519);
    sample_manager_inst.add_one_monitor(fifo_monitor_520);
    sample_manager_inst.add_one_monitor(fifo_monitor_521);
    sample_manager_inst.add_one_monitor(fifo_monitor_522);
    sample_manager_inst.add_one_monitor(fifo_monitor_523);
    sample_manager_inst.add_one_monitor(fifo_monitor_524);
    sample_manager_inst.add_one_monitor(fifo_monitor_525);
    sample_manager_inst.add_one_monitor(fifo_monitor_526);
    sample_manager_inst.add_one_monitor(fifo_monitor_527);
    sample_manager_inst.add_one_monitor(fifo_monitor_528);
    sample_manager_inst.add_one_monitor(fifo_monitor_529);
    sample_manager_inst.add_one_monitor(fifo_monitor_530);
    sample_manager_inst.add_one_monitor(fifo_monitor_531);
    sample_manager_inst.add_one_monitor(fifo_monitor_532);
    sample_manager_inst.add_one_monitor(fifo_monitor_533);
    sample_manager_inst.add_one_monitor(fifo_monitor_534);
    sample_manager_inst.add_one_monitor(fifo_monitor_535);
    sample_manager_inst.add_one_monitor(fifo_monitor_536);
    sample_manager_inst.add_one_monitor(fifo_monitor_537);
    sample_manager_inst.add_one_monitor(fifo_monitor_538);
    sample_manager_inst.add_one_monitor(fifo_monitor_539);
    sample_manager_inst.add_one_monitor(fifo_monitor_540);
    sample_manager_inst.add_one_monitor(fifo_monitor_541);
    sample_manager_inst.add_one_monitor(fifo_monitor_542);
    sample_manager_inst.add_one_monitor(fifo_monitor_543);
    sample_manager_inst.add_one_monitor(fifo_monitor_544);
    sample_manager_inst.add_one_monitor(fifo_monitor_545);
    sample_manager_inst.add_one_monitor(fifo_monitor_546);
    sample_manager_inst.add_one_monitor(fifo_monitor_547);
    sample_manager_inst.add_one_monitor(fifo_monitor_548);
    sample_manager_inst.add_one_monitor(fifo_monitor_549);
    sample_manager_inst.add_one_monitor(fifo_monitor_550);
    sample_manager_inst.add_one_monitor(fifo_monitor_551);
    sample_manager_inst.add_one_monitor(fifo_monitor_552);
    sample_manager_inst.add_one_monitor(fifo_monitor_553);
    sample_manager_inst.add_one_monitor(fifo_monitor_554);
    sample_manager_inst.add_one_monitor(fifo_monitor_555);
    sample_manager_inst.add_one_monitor(fifo_monitor_556);
    sample_manager_inst.add_one_monitor(fifo_monitor_557);
    sample_manager_inst.add_one_monitor(fifo_monitor_558);
    sample_manager_inst.add_one_monitor(fifo_monitor_559);
    sample_manager_inst.add_one_monitor(fifo_monitor_560);
    sample_manager_inst.add_one_monitor(fifo_monitor_561);
    sample_manager_inst.add_one_monitor(fifo_monitor_562);
    sample_manager_inst.add_one_monitor(fifo_monitor_563);
    sample_manager_inst.add_one_monitor(fifo_monitor_564);
    sample_manager_inst.add_one_monitor(fifo_monitor_565);
    sample_manager_inst.add_one_monitor(fifo_monitor_566);
    sample_manager_inst.add_one_monitor(fifo_monitor_567);
    sample_manager_inst.add_one_monitor(fifo_monitor_568);
    sample_manager_inst.add_one_monitor(fifo_monitor_569);
    sample_manager_inst.add_one_monitor(fifo_monitor_570);
    sample_manager_inst.add_one_monitor(fifo_monitor_571);
    sample_manager_inst.add_one_monitor(fifo_monitor_572);
    sample_manager_inst.add_one_monitor(fifo_monitor_573);
    sample_manager_inst.add_one_monitor(fifo_monitor_574);
    sample_manager_inst.add_one_monitor(fifo_monitor_575);
    sample_manager_inst.add_one_monitor(fifo_monitor_576);
    sample_manager_inst.add_one_monitor(fifo_monitor_577);
    sample_manager_inst.add_one_monitor(fifo_monitor_578);
    sample_manager_inst.add_one_monitor(fifo_monitor_579);
    sample_manager_inst.add_one_monitor(fifo_monitor_580);
    sample_manager_inst.add_one_monitor(fifo_monitor_581);
    sample_manager_inst.add_one_monitor(fifo_monitor_582);
    sample_manager_inst.add_one_monitor(fifo_monitor_583);
    sample_manager_inst.add_one_monitor(fifo_monitor_584);
    sample_manager_inst.add_one_monitor(fifo_monitor_585);
    sample_manager_inst.add_one_monitor(fifo_monitor_586);
    sample_manager_inst.add_one_monitor(fifo_monitor_587);
    sample_manager_inst.add_one_monitor(fifo_monitor_588);
    sample_manager_inst.add_one_monitor(fifo_monitor_589);
    sample_manager_inst.add_one_monitor(fifo_monitor_590);
    sample_manager_inst.add_one_monitor(fifo_monitor_591);
    sample_manager_inst.add_one_monitor(fifo_monitor_592);
    sample_manager_inst.add_one_monitor(fifo_monitor_593);
    sample_manager_inst.add_one_monitor(fifo_monitor_594);
    sample_manager_inst.add_one_monitor(fifo_monitor_595);
    sample_manager_inst.add_one_monitor(fifo_monitor_596);
    sample_manager_inst.add_one_monitor(fifo_monitor_597);
    sample_manager_inst.add_one_monitor(fifo_monitor_598);
    sample_manager_inst.add_one_monitor(fifo_monitor_599);
    sample_manager_inst.add_one_monitor(fifo_monitor_600);
    sample_manager_inst.add_one_monitor(fifo_monitor_601);
    sample_manager_inst.add_one_monitor(fifo_monitor_602);
    sample_manager_inst.add_one_monitor(fifo_monitor_603);
    sample_manager_inst.add_one_monitor(fifo_monitor_604);
    sample_manager_inst.add_one_monitor(fifo_monitor_605);
    sample_manager_inst.add_one_monitor(fifo_monitor_606);
    sample_manager_inst.add_one_monitor(fifo_monitor_607);
    sample_manager_inst.add_one_monitor(fifo_monitor_608);
    sample_manager_inst.add_one_monitor(fifo_monitor_609);
    sample_manager_inst.add_one_monitor(fifo_monitor_610);
    sample_manager_inst.add_one_monitor(fifo_monitor_611);
    sample_manager_inst.add_one_monitor(fifo_monitor_612);
    sample_manager_inst.add_one_monitor(fifo_monitor_613);
    sample_manager_inst.add_one_monitor(fifo_monitor_614);
    sample_manager_inst.add_one_monitor(fifo_monitor_615);
    sample_manager_inst.add_one_monitor(fifo_monitor_616);
    sample_manager_inst.add_one_monitor(fifo_monitor_617);
    sample_manager_inst.add_one_monitor(fifo_monitor_618);
    sample_manager_inst.add_one_monitor(fifo_monitor_619);
    sample_manager_inst.add_one_monitor(fifo_monitor_620);
    sample_manager_inst.add_one_monitor(fifo_monitor_621);
    sample_manager_inst.add_one_monitor(fifo_monitor_622);
    sample_manager_inst.add_one_monitor(fifo_monitor_623);
    sample_manager_inst.add_one_monitor(fifo_monitor_624);
    sample_manager_inst.add_one_monitor(fifo_monitor_625);
    sample_manager_inst.add_one_monitor(fifo_monitor_626);
    sample_manager_inst.add_one_monitor(fifo_monitor_627);
    sample_manager_inst.add_one_monitor(fifo_monitor_628);
    sample_manager_inst.add_one_monitor(fifo_monitor_629);
    sample_manager_inst.add_one_monitor(fifo_monitor_630);
    sample_manager_inst.add_one_monitor(fifo_monitor_631);
    sample_manager_inst.add_one_monitor(fifo_monitor_632);
    sample_manager_inst.add_one_monitor(fifo_monitor_633);
    sample_manager_inst.add_one_monitor(fifo_monitor_634);
    sample_manager_inst.add_one_monitor(fifo_monitor_635);
    sample_manager_inst.add_one_monitor(fifo_monitor_636);
    sample_manager_inst.add_one_monitor(fifo_monitor_637);
    sample_manager_inst.add_one_monitor(fifo_monitor_638);
    sample_manager_inst.add_one_monitor(fifo_monitor_639);
    sample_manager_inst.add_one_monitor(fifo_monitor_640);
    sample_manager_inst.add_one_monitor(fifo_monitor_641);
    sample_manager_inst.add_one_monitor(fifo_monitor_642);
    sample_manager_inst.add_one_monitor(fifo_monitor_643);
    sample_manager_inst.add_one_monitor(fifo_monitor_644);
    sample_manager_inst.add_one_monitor(fifo_monitor_645);
    sample_manager_inst.add_one_monitor(fifo_monitor_646);
    sample_manager_inst.add_one_monitor(fifo_monitor_647);
    sample_manager_inst.add_one_monitor(fifo_monitor_648);
    sample_manager_inst.add_one_monitor(fifo_monitor_649);
    sample_manager_inst.add_one_monitor(fifo_monitor_650);
    sample_manager_inst.add_one_monitor(fifo_monitor_651);
    sample_manager_inst.add_one_monitor(fifo_monitor_652);
    sample_manager_inst.add_one_monitor(fifo_monitor_653);
    sample_manager_inst.add_one_monitor(fifo_monitor_654);
    sample_manager_inst.add_one_monitor(fifo_monitor_655);
    sample_manager_inst.add_one_monitor(fifo_monitor_656);
    sample_manager_inst.add_one_monitor(fifo_monitor_657);
    sample_manager_inst.add_one_monitor(fifo_monitor_658);
    sample_manager_inst.add_one_monitor(fifo_monitor_659);
    sample_manager_inst.add_one_monitor(fifo_monitor_660);
    sample_manager_inst.add_one_monitor(fifo_monitor_661);
    sample_manager_inst.add_one_monitor(fifo_monitor_662);
    sample_manager_inst.add_one_monitor(fifo_monitor_663);
    sample_manager_inst.add_one_monitor(fifo_monitor_664);
    sample_manager_inst.add_one_monitor(fifo_monitor_665);
    sample_manager_inst.add_one_monitor(fifo_monitor_666);
    sample_manager_inst.add_one_monitor(fifo_monitor_667);
    sample_manager_inst.add_one_monitor(fifo_monitor_668);
    sample_manager_inst.add_one_monitor(fifo_monitor_669);
    sample_manager_inst.add_one_monitor(fifo_monitor_670);
    sample_manager_inst.add_one_monitor(fifo_monitor_671);
    sample_manager_inst.add_one_monitor(fifo_monitor_672);
    sample_manager_inst.add_one_monitor(fifo_monitor_673);
    sample_manager_inst.add_one_monitor(fifo_monitor_674);
    sample_manager_inst.add_one_monitor(fifo_monitor_675);
    sample_manager_inst.add_one_monitor(fifo_monitor_676);
    sample_manager_inst.add_one_monitor(fifo_monitor_677);
    sample_manager_inst.add_one_monitor(fifo_monitor_678);
    sample_manager_inst.add_one_monitor(fifo_monitor_679);
    sample_manager_inst.add_one_monitor(fifo_monitor_680);
    sample_manager_inst.add_one_monitor(fifo_monitor_681);
    sample_manager_inst.add_one_monitor(fifo_monitor_682);
    sample_manager_inst.add_one_monitor(fifo_monitor_683);
    sample_manager_inst.add_one_monitor(fifo_monitor_684);
    sample_manager_inst.add_one_monitor(fifo_monitor_685);
    sample_manager_inst.add_one_monitor(fifo_monitor_686);
    sample_manager_inst.add_one_monitor(fifo_monitor_687);
    sample_manager_inst.add_one_monitor(fifo_monitor_688);
    sample_manager_inst.add_one_monitor(fifo_monitor_689);
    sample_manager_inst.add_one_monitor(fifo_monitor_690);
    sample_manager_inst.add_one_monitor(fifo_monitor_691);
    sample_manager_inst.add_one_monitor(fifo_monitor_692);
    sample_manager_inst.add_one_monitor(fifo_monitor_693);
    sample_manager_inst.add_one_monitor(fifo_monitor_694);
    sample_manager_inst.add_one_monitor(fifo_monitor_695);
    sample_manager_inst.add_one_monitor(fifo_monitor_696);
    sample_manager_inst.add_one_monitor(fifo_monitor_697);
    sample_manager_inst.add_one_monitor(fifo_monitor_698);
    sample_manager_inst.add_one_monitor(fifo_monitor_699);
    sample_manager_inst.add_one_monitor(fifo_monitor_700);
    sample_manager_inst.add_one_monitor(fifo_monitor_701);
    sample_manager_inst.add_one_monitor(fifo_monitor_702);
    sample_manager_inst.add_one_monitor(fifo_monitor_703);
    sample_manager_inst.add_one_monitor(fifo_monitor_704);
    sample_manager_inst.add_one_monitor(fifo_monitor_705);
    sample_manager_inst.add_one_monitor(fifo_monitor_706);
    sample_manager_inst.add_one_monitor(fifo_monitor_707);
    sample_manager_inst.add_one_monitor(fifo_monitor_708);
    sample_manager_inst.add_one_monitor(fifo_monitor_709);
    sample_manager_inst.add_one_monitor(fifo_monitor_710);
    sample_manager_inst.add_one_monitor(fifo_monitor_711);
    sample_manager_inst.add_one_monitor(fifo_monitor_712);
    sample_manager_inst.add_one_monitor(fifo_monitor_713);
    sample_manager_inst.add_one_monitor(fifo_monitor_714);
    sample_manager_inst.add_one_monitor(fifo_monitor_715);
    sample_manager_inst.add_one_monitor(fifo_monitor_716);
    sample_manager_inst.add_one_monitor(fifo_monitor_717);
    sample_manager_inst.add_one_monitor(fifo_monitor_718);
    sample_manager_inst.add_one_monitor(fifo_monitor_719);
    sample_manager_inst.add_one_monitor(fifo_monitor_720);
    sample_manager_inst.add_one_monitor(fifo_monitor_721);
    sample_manager_inst.add_one_monitor(fifo_monitor_722);
    sample_manager_inst.add_one_monitor(fifo_monitor_723);
    sample_manager_inst.add_one_monitor(fifo_monitor_724);
    sample_manager_inst.add_one_monitor(fifo_monitor_725);
    sample_manager_inst.add_one_monitor(fifo_monitor_726);
    sample_manager_inst.add_one_monitor(fifo_monitor_727);
    sample_manager_inst.add_one_monitor(fifo_monitor_728);
    sample_manager_inst.add_one_monitor(fifo_monitor_729);
    sample_manager_inst.add_one_monitor(fifo_monitor_730);
    sample_manager_inst.add_one_monitor(fifo_monitor_731);
    sample_manager_inst.add_one_monitor(fifo_monitor_732);
    sample_manager_inst.add_one_monitor(fifo_monitor_733);
    sample_manager_inst.add_one_monitor(fifo_monitor_734);
    sample_manager_inst.add_one_monitor(fifo_monitor_735);
    sample_manager_inst.add_one_monitor(fifo_monitor_736);
    sample_manager_inst.add_one_monitor(fifo_monitor_737);
    sample_manager_inst.add_one_monitor(fifo_monitor_738);
    sample_manager_inst.add_one_monitor(fifo_monitor_739);
    sample_manager_inst.add_one_monitor(fifo_monitor_740);
    sample_manager_inst.add_one_monitor(fifo_monitor_741);
    sample_manager_inst.add_one_monitor(fifo_monitor_742);
    sample_manager_inst.add_one_monitor(fifo_monitor_743);
    sample_manager_inst.add_one_monitor(fifo_monitor_744);
    sample_manager_inst.add_one_monitor(fifo_monitor_745);
    sample_manager_inst.add_one_monitor(fifo_monitor_746);
    sample_manager_inst.add_one_monitor(fifo_monitor_747);
    sample_manager_inst.add_one_monitor(fifo_monitor_748);
    sample_manager_inst.add_one_monitor(fifo_monitor_749);
    sample_manager_inst.add_one_monitor(fifo_monitor_750);
    sample_manager_inst.add_one_monitor(fifo_monitor_751);
    sample_manager_inst.add_one_monitor(fifo_monitor_752);
    sample_manager_inst.add_one_monitor(fifo_monitor_753);
    sample_manager_inst.add_one_monitor(fifo_monitor_754);
    sample_manager_inst.add_one_monitor(fifo_monitor_755);
    sample_manager_inst.add_one_monitor(fifo_monitor_756);
    sample_manager_inst.add_one_monitor(fifo_monitor_757);
    sample_manager_inst.add_one_monitor(fifo_monitor_758);
    sample_manager_inst.add_one_monitor(fifo_monitor_759);
    sample_manager_inst.add_one_monitor(fifo_monitor_760);
    sample_manager_inst.add_one_monitor(fifo_monitor_761);
    sample_manager_inst.add_one_monitor(fifo_monitor_762);
    sample_manager_inst.add_one_monitor(fifo_monitor_763);
    sample_manager_inst.add_one_monitor(fifo_monitor_764);
    sample_manager_inst.add_one_monitor(fifo_monitor_765);
    sample_manager_inst.add_one_monitor(fifo_monitor_766);
    sample_manager_inst.add_one_monitor(fifo_monitor_767);
    sample_manager_inst.add_one_monitor(fifo_monitor_768);
    sample_manager_inst.add_one_monitor(fifo_monitor_769);
    sample_manager_inst.add_one_monitor(fifo_monitor_770);
    sample_manager_inst.add_one_monitor(fifo_monitor_771);
    sample_manager_inst.add_one_monitor(fifo_monitor_772);
    sample_manager_inst.add_one_monitor(fifo_monitor_773);
    sample_manager_inst.add_one_monitor(fifo_monitor_774);
    sample_manager_inst.add_one_monitor(fifo_monitor_775);
    sample_manager_inst.add_one_monitor(fifo_monitor_776);
    sample_manager_inst.add_one_monitor(fifo_monitor_777);
    sample_manager_inst.add_one_monitor(fifo_monitor_778);
    sample_manager_inst.add_one_monitor(fifo_monitor_779);
    sample_manager_inst.add_one_monitor(fifo_monitor_780);
    sample_manager_inst.add_one_monitor(fifo_monitor_781);
    sample_manager_inst.add_one_monitor(fifo_monitor_782);
    sample_manager_inst.add_one_monitor(fifo_monitor_783);
    sample_manager_inst.add_one_monitor(fifo_monitor_784);
    sample_manager_inst.add_one_monitor(fifo_monitor_785);
    sample_manager_inst.add_one_monitor(fifo_monitor_786);
    sample_manager_inst.add_one_monitor(fifo_monitor_787);
    sample_manager_inst.add_one_monitor(fifo_monitor_788);
    sample_manager_inst.add_one_monitor(fifo_monitor_789);
    sample_manager_inst.add_one_monitor(fifo_monitor_790);
    sample_manager_inst.add_one_monitor(fifo_monitor_791);
    sample_manager_inst.add_one_monitor(fifo_monitor_792);
    sample_manager_inst.add_one_monitor(fifo_monitor_793);
    sample_manager_inst.add_one_monitor(fifo_monitor_794);
    sample_manager_inst.add_one_monitor(fifo_monitor_795);
    sample_manager_inst.add_one_monitor(fifo_monitor_796);
    sample_manager_inst.add_one_monitor(fifo_monitor_797);
    sample_manager_inst.add_one_monitor(fifo_monitor_798);
    sample_manager_inst.add_one_monitor(fifo_monitor_799);
    sample_manager_inst.add_one_monitor(fifo_monitor_800);
    sample_manager_inst.add_one_monitor(fifo_monitor_801);
    sample_manager_inst.add_one_monitor(fifo_monitor_802);
    sample_manager_inst.add_one_monitor(fifo_monitor_803);
    sample_manager_inst.add_one_monitor(fifo_monitor_804);
    sample_manager_inst.add_one_monitor(fifo_monitor_805);
    sample_manager_inst.add_one_monitor(fifo_monitor_806);
    sample_manager_inst.add_one_monitor(fifo_monitor_807);
    sample_manager_inst.add_one_monitor(fifo_monitor_808);
    sample_manager_inst.add_one_monitor(fifo_monitor_809);
    sample_manager_inst.add_one_monitor(fifo_monitor_810);
    sample_manager_inst.add_one_monitor(fifo_monitor_811);
    sample_manager_inst.add_one_monitor(fifo_monitor_812);
    sample_manager_inst.add_one_monitor(fifo_monitor_813);
    sample_manager_inst.add_one_monitor(fifo_monitor_814);
    sample_manager_inst.add_one_monitor(fifo_monitor_815);
    sample_manager_inst.add_one_monitor(fifo_monitor_816);
    sample_manager_inst.add_one_monitor(fifo_monitor_817);
    sample_manager_inst.add_one_monitor(fifo_monitor_818);
    sample_manager_inst.add_one_monitor(fifo_monitor_819);
    sample_manager_inst.add_one_monitor(fifo_monitor_820);
    sample_manager_inst.add_one_monitor(fifo_monitor_821);
    sample_manager_inst.add_one_monitor(fifo_monitor_822);
    sample_manager_inst.add_one_monitor(fifo_monitor_823);
    sample_manager_inst.add_one_monitor(fifo_monitor_824);
    sample_manager_inst.add_one_monitor(fifo_monitor_825);
    sample_manager_inst.add_one_monitor(fifo_monitor_826);
    sample_manager_inst.add_one_monitor(fifo_monitor_827);
    sample_manager_inst.add_one_monitor(fifo_monitor_828);
    sample_manager_inst.add_one_monitor(fifo_monitor_829);
    sample_manager_inst.add_one_monitor(fifo_monitor_830);
    sample_manager_inst.add_one_monitor(fifo_monitor_831);
    sample_manager_inst.add_one_monitor(fifo_monitor_832);
    sample_manager_inst.add_one_monitor(fifo_monitor_833);
    sample_manager_inst.add_one_monitor(fifo_monitor_834);
    sample_manager_inst.add_one_monitor(fifo_monitor_835);
    sample_manager_inst.add_one_monitor(fifo_monitor_836);
    sample_manager_inst.add_one_monitor(fifo_monitor_837);
    sample_manager_inst.add_one_monitor(fifo_monitor_838);
    sample_manager_inst.add_one_monitor(fifo_monitor_839);
    sample_manager_inst.add_one_monitor(fifo_monitor_840);
    sample_manager_inst.add_one_monitor(fifo_monitor_841);
    sample_manager_inst.add_one_monitor(fifo_monitor_842);
    sample_manager_inst.add_one_monitor(fifo_monitor_843);
    sample_manager_inst.add_one_monitor(fifo_monitor_844);
    sample_manager_inst.add_one_monitor(fifo_monitor_845);
    sample_manager_inst.add_one_monitor(fifo_monitor_846);
    sample_manager_inst.add_one_monitor(fifo_monitor_847);
    sample_manager_inst.add_one_monitor(fifo_monitor_848);
    sample_manager_inst.add_one_monitor(fifo_monitor_849);
    sample_manager_inst.add_one_monitor(fifo_monitor_850);
    sample_manager_inst.add_one_monitor(fifo_monitor_851);
    sample_manager_inst.add_one_monitor(fifo_monitor_852);
    sample_manager_inst.add_one_monitor(fifo_monitor_853);
    sample_manager_inst.add_one_monitor(fifo_monitor_854);
    sample_manager_inst.add_one_monitor(fifo_monitor_855);
    sample_manager_inst.add_one_monitor(fifo_monitor_856);
    sample_manager_inst.add_one_monitor(fifo_monitor_857);
    sample_manager_inst.add_one_monitor(fifo_monitor_858);
    sample_manager_inst.add_one_monitor(fifo_monitor_859);
    sample_manager_inst.add_one_monitor(fifo_monitor_860);
    sample_manager_inst.add_one_monitor(fifo_monitor_861);
    sample_manager_inst.add_one_monitor(fifo_monitor_862);
    sample_manager_inst.add_one_monitor(fifo_monitor_863);
    sample_manager_inst.add_one_monitor(fifo_monitor_864);
    sample_manager_inst.add_one_monitor(fifo_monitor_865);
    sample_manager_inst.add_one_monitor(fifo_monitor_866);
    sample_manager_inst.add_one_monitor(fifo_monitor_867);
    sample_manager_inst.add_one_monitor(fifo_monitor_868);
    sample_manager_inst.add_one_monitor(fifo_monitor_869);
    sample_manager_inst.add_one_monitor(fifo_monitor_870);
    sample_manager_inst.add_one_monitor(fifo_monitor_871);
    sample_manager_inst.add_one_monitor(fifo_monitor_872);
    sample_manager_inst.add_one_monitor(fifo_monitor_873);
    sample_manager_inst.add_one_monitor(fifo_monitor_874);
    sample_manager_inst.add_one_monitor(fifo_monitor_875);
    sample_manager_inst.add_one_monitor(fifo_monitor_876);
    sample_manager_inst.add_one_monitor(fifo_monitor_877);
    sample_manager_inst.add_one_monitor(fifo_monitor_878);
    sample_manager_inst.add_one_monitor(fifo_monitor_879);
    sample_manager_inst.add_one_monitor(fifo_monitor_880);
    sample_manager_inst.add_one_monitor(fifo_monitor_881);
    sample_manager_inst.add_one_monitor(fifo_monitor_882);
    sample_manager_inst.add_one_monitor(fifo_monitor_883);
    sample_manager_inst.add_one_monitor(fifo_monitor_884);
    sample_manager_inst.add_one_monitor(fifo_monitor_885);
    sample_manager_inst.add_one_monitor(fifo_monitor_886);
    sample_manager_inst.add_one_monitor(fifo_monitor_887);
    sample_manager_inst.add_one_monitor(fifo_monitor_888);
    sample_manager_inst.add_one_monitor(fifo_monitor_889);
    sample_manager_inst.add_one_monitor(fifo_monitor_890);
    sample_manager_inst.add_one_monitor(fifo_monitor_891);
    sample_manager_inst.add_one_monitor(fifo_monitor_892);
    sample_manager_inst.add_one_monitor(fifo_monitor_893);
    sample_manager_inst.add_one_monitor(fifo_monitor_894);
    sample_manager_inst.add_one_monitor(fifo_monitor_895);
    sample_manager_inst.add_one_monitor(fifo_monitor_896);
    sample_manager_inst.add_one_monitor(fifo_monitor_897);
    sample_manager_inst.add_one_monitor(fifo_monitor_898);
    sample_manager_inst.add_one_monitor(fifo_monitor_899);
    sample_manager_inst.add_one_monitor(fifo_monitor_900);
    sample_manager_inst.add_one_monitor(fifo_monitor_901);
    sample_manager_inst.add_one_monitor(fifo_monitor_902);
    sample_manager_inst.add_one_monitor(fifo_monitor_903);
    sample_manager_inst.add_one_monitor(fifo_monitor_904);
    sample_manager_inst.add_one_monitor(fifo_monitor_905);
    sample_manager_inst.add_one_monitor(fifo_monitor_906);
    sample_manager_inst.add_one_monitor(fifo_monitor_907);
    sample_manager_inst.add_one_monitor(fifo_monitor_908);
    sample_manager_inst.add_one_monitor(fifo_monitor_909);
    sample_manager_inst.add_one_monitor(fifo_monitor_910);
    sample_manager_inst.add_one_monitor(fifo_monitor_911);
    sample_manager_inst.add_one_monitor(fifo_monitor_912);
    sample_manager_inst.add_one_monitor(fifo_monitor_913);
    sample_manager_inst.add_one_monitor(fifo_monitor_914);
    sample_manager_inst.add_one_monitor(fifo_monitor_915);
    sample_manager_inst.add_one_monitor(fifo_monitor_916);
    sample_manager_inst.add_one_monitor(fifo_monitor_917);
    sample_manager_inst.add_one_monitor(fifo_monitor_918);
    sample_manager_inst.add_one_monitor(fifo_monitor_919);
    sample_manager_inst.add_one_monitor(fifo_monitor_920);
    sample_manager_inst.add_one_monitor(fifo_monitor_921);
    sample_manager_inst.add_one_monitor(fifo_monitor_922);
    sample_manager_inst.add_one_monitor(fifo_monitor_923);
    sample_manager_inst.add_one_monitor(fifo_monitor_924);
    sample_manager_inst.add_one_monitor(fifo_monitor_925);
    sample_manager_inst.add_one_monitor(fifo_monitor_926);
    sample_manager_inst.add_one_monitor(fifo_monitor_927);
    sample_manager_inst.add_one_monitor(fifo_monitor_928);
    sample_manager_inst.add_one_monitor(fifo_monitor_929);
    sample_manager_inst.add_one_monitor(fifo_monitor_930);
    sample_manager_inst.add_one_monitor(fifo_monitor_931);
    sample_manager_inst.add_one_monitor(fifo_monitor_932);
    sample_manager_inst.add_one_monitor(fifo_monitor_933);
    sample_manager_inst.add_one_monitor(fifo_monitor_934);
    sample_manager_inst.add_one_monitor(fifo_monitor_935);
    sample_manager_inst.add_one_monitor(fifo_monitor_936);
    sample_manager_inst.add_one_monitor(fifo_monitor_937);
    sample_manager_inst.add_one_monitor(fifo_monitor_938);
    sample_manager_inst.add_one_monitor(fifo_monitor_939);
    sample_manager_inst.add_one_monitor(fifo_monitor_940);
    sample_manager_inst.add_one_monitor(fifo_monitor_941);
    sample_manager_inst.add_one_monitor(fifo_monitor_942);
    sample_manager_inst.add_one_monitor(fifo_monitor_943);
    sample_manager_inst.add_one_monitor(fifo_monitor_944);
    sample_manager_inst.add_one_monitor(fifo_monitor_945);
    sample_manager_inst.add_one_monitor(fifo_monitor_946);
    sample_manager_inst.add_one_monitor(fifo_monitor_947);
    sample_manager_inst.add_one_monitor(fifo_monitor_948);
    sample_manager_inst.add_one_monitor(fifo_monitor_949);
    sample_manager_inst.add_one_monitor(fifo_monitor_950);
    sample_manager_inst.add_one_monitor(fifo_monitor_951);
    sample_manager_inst.add_one_monitor(fifo_monitor_952);
    sample_manager_inst.add_one_monitor(fifo_monitor_953);
    sample_manager_inst.add_one_monitor(fifo_monitor_954);
    sample_manager_inst.add_one_monitor(fifo_monitor_955);
    sample_manager_inst.add_one_monitor(fifo_monitor_956);
    sample_manager_inst.add_one_monitor(fifo_monitor_957);
    sample_manager_inst.add_one_monitor(fifo_monitor_958);
    sample_manager_inst.add_one_monitor(fifo_monitor_959);
    sample_manager_inst.add_one_monitor(fifo_monitor_960);
    sample_manager_inst.add_one_monitor(fifo_monitor_961);
    sample_manager_inst.add_one_monitor(fifo_monitor_962);
    sample_manager_inst.add_one_monitor(fifo_monitor_963);
    sample_manager_inst.add_one_monitor(fifo_monitor_964);
    sample_manager_inst.add_one_monitor(fifo_monitor_965);
    sample_manager_inst.add_one_monitor(fifo_monitor_966);
    sample_manager_inst.add_one_monitor(fifo_monitor_967);
    sample_manager_inst.add_one_monitor(fifo_monitor_968);
    sample_manager_inst.add_one_monitor(fifo_monitor_969);
    sample_manager_inst.add_one_monitor(fifo_monitor_970);
    sample_manager_inst.add_one_monitor(fifo_monitor_971);
    sample_manager_inst.add_one_monitor(fifo_monitor_972);
    sample_manager_inst.add_one_monitor(fifo_monitor_973);
    sample_manager_inst.add_one_monitor(fifo_monitor_974);
    sample_manager_inst.add_one_monitor(fifo_monitor_975);
    sample_manager_inst.add_one_monitor(fifo_monitor_976);
    sample_manager_inst.add_one_monitor(fifo_monitor_977);
    sample_manager_inst.add_one_monitor(fifo_monitor_978);
    sample_manager_inst.add_one_monitor(fifo_monitor_979);
    sample_manager_inst.add_one_monitor(fifo_monitor_980);
    sample_manager_inst.add_one_monitor(fifo_monitor_981);
    sample_manager_inst.add_one_monitor(fifo_monitor_982);
    sample_manager_inst.add_one_monitor(fifo_monitor_983);
    sample_manager_inst.add_one_monitor(fifo_monitor_984);
    sample_manager_inst.add_one_monitor(fifo_monitor_985);
    sample_manager_inst.add_one_monitor(fifo_monitor_986);
    sample_manager_inst.add_one_monitor(fifo_monitor_987);
    sample_manager_inst.add_one_monitor(fifo_monitor_988);
    sample_manager_inst.add_one_monitor(fifo_monitor_989);
    sample_manager_inst.add_one_monitor(fifo_monitor_990);
    sample_manager_inst.add_one_monitor(fifo_monitor_991);
    sample_manager_inst.add_one_monitor(fifo_monitor_992);
    sample_manager_inst.add_one_monitor(fifo_monitor_993);
    sample_manager_inst.add_one_monitor(fifo_monitor_994);
    sample_manager_inst.add_one_monitor(fifo_monitor_995);
    sample_manager_inst.add_one_monitor(fifo_monitor_996);
    sample_manager_inst.add_one_monitor(fifo_monitor_997);
    sample_manager_inst.add_one_monitor(fifo_monitor_998);
    sample_manager_inst.add_one_monitor(fifo_monitor_999);
    sample_manager_inst.add_one_monitor(fifo_monitor_1000);
    sample_manager_inst.add_one_monitor(fifo_monitor_1001);
    sample_manager_inst.add_one_monitor(fifo_monitor_1002);
    sample_manager_inst.add_one_monitor(fifo_monitor_1003);
    sample_manager_inst.add_one_monitor(fifo_monitor_1004);
    sample_manager_inst.add_one_monitor(fifo_monitor_1005);
    sample_manager_inst.add_one_monitor(fifo_monitor_1006);
    sample_manager_inst.add_one_monitor(fifo_monitor_1007);
    sample_manager_inst.add_one_monitor(fifo_monitor_1008);
    sample_manager_inst.add_one_monitor(fifo_monitor_1009);
    sample_manager_inst.add_one_monitor(fifo_monitor_1010);
    sample_manager_inst.add_one_monitor(fifo_monitor_1011);
    sample_manager_inst.add_one_monitor(fifo_monitor_1012);
    sample_manager_inst.add_one_monitor(fifo_monitor_1013);
    sample_manager_inst.add_one_monitor(fifo_monitor_1014);
    sample_manager_inst.add_one_monitor(fifo_monitor_1015);
    sample_manager_inst.add_one_monitor(fifo_monitor_1016);
    sample_manager_inst.add_one_monitor(fifo_monitor_1017);
    sample_manager_inst.add_one_monitor(fifo_monitor_1018);
    sample_manager_inst.add_one_monitor(fifo_monitor_1019);
    sample_manager_inst.add_one_monitor(fifo_monitor_1020);
    sample_manager_inst.add_one_monitor(fifo_monitor_1021);
    sample_manager_inst.add_one_monitor(fifo_monitor_1022);
    sample_manager_inst.add_one_monitor(fifo_monitor_1023);
    sample_manager_inst.add_one_monitor(fifo_monitor_1024);
    sample_manager_inst.add_one_monitor(fifo_monitor_1025);
    sample_manager_inst.add_one_monitor(fifo_monitor_1026);
    sample_manager_inst.add_one_monitor(fifo_monitor_1027);
    sample_manager_inst.add_one_monitor(fifo_monitor_1028);
    sample_manager_inst.add_one_monitor(fifo_monitor_1029);
    sample_manager_inst.add_one_monitor(fifo_monitor_1030);
    sample_manager_inst.add_one_monitor(fifo_monitor_1031);
    sample_manager_inst.add_one_monitor(fifo_monitor_1032);
    sample_manager_inst.add_one_monitor(fifo_monitor_1033);
    sample_manager_inst.add_one_monitor(fifo_monitor_1034);
    sample_manager_inst.add_one_monitor(fifo_monitor_1035);
    sample_manager_inst.add_one_monitor(fifo_monitor_1036);
    sample_manager_inst.add_one_monitor(fifo_monitor_1037);
    sample_manager_inst.add_one_monitor(fifo_monitor_1038);
    sample_manager_inst.add_one_monitor(fifo_monitor_1039);
    sample_manager_inst.add_one_monitor(fifo_monitor_1040);
    sample_manager_inst.add_one_monitor(fifo_monitor_1041);
    sample_manager_inst.add_one_monitor(fifo_monitor_1042);
    sample_manager_inst.add_one_monitor(fifo_monitor_1043);
    sample_manager_inst.add_one_monitor(fifo_monitor_1044);
    sample_manager_inst.add_one_monitor(fifo_monitor_1045);
    sample_manager_inst.add_one_monitor(fifo_monitor_1046);
    sample_manager_inst.add_one_monitor(fifo_monitor_1047);
    sample_manager_inst.add_one_monitor(fifo_monitor_1048);
    sample_manager_inst.add_one_monitor(fifo_monitor_1049);
    sample_manager_inst.add_one_monitor(fifo_monitor_1050);
    sample_manager_inst.add_one_monitor(fifo_monitor_1051);
    sample_manager_inst.add_one_monitor(fifo_monitor_1052);
    sample_manager_inst.add_one_monitor(fifo_monitor_1053);
    sample_manager_inst.add_one_monitor(fifo_monitor_1054);
    sample_manager_inst.add_one_monitor(fifo_monitor_1055);
    sample_manager_inst.add_one_monitor(fifo_monitor_1056);
    sample_manager_inst.add_one_monitor(fifo_monitor_1057);
    sample_manager_inst.add_one_monitor(fifo_monitor_1058);
    sample_manager_inst.add_one_monitor(fifo_monitor_1059);
    sample_manager_inst.add_one_monitor(fifo_monitor_1060);
    sample_manager_inst.add_one_monitor(fifo_monitor_1061);
    sample_manager_inst.add_one_monitor(fifo_monitor_1062);
    sample_manager_inst.add_one_monitor(fifo_monitor_1063);
    sample_manager_inst.add_one_monitor(fifo_monitor_1064);
    sample_manager_inst.add_one_monitor(fifo_monitor_1065);
    sample_manager_inst.add_one_monitor(fifo_monitor_1066);
    sample_manager_inst.add_one_monitor(fifo_monitor_1067);
    sample_manager_inst.add_one_monitor(fifo_monitor_1068);
    sample_manager_inst.add_one_monitor(fifo_monitor_1069);
    sample_manager_inst.add_one_monitor(fifo_monitor_1070);
    sample_manager_inst.add_one_monitor(fifo_monitor_1071);
    sample_manager_inst.add_one_monitor(fifo_monitor_1072);
    sample_manager_inst.add_one_monitor(fifo_monitor_1073);
    sample_manager_inst.add_one_monitor(fifo_monitor_1074);
    sample_manager_inst.add_one_monitor(fifo_monitor_1075);
    sample_manager_inst.add_one_monitor(fifo_monitor_1076);
    sample_manager_inst.add_one_monitor(fifo_monitor_1077);
    sample_manager_inst.add_one_monitor(fifo_monitor_1078);
    sample_manager_inst.add_one_monitor(fifo_monitor_1079);
    sample_manager_inst.add_one_monitor(fifo_monitor_1080);
    sample_manager_inst.add_one_monitor(fifo_monitor_1081);
    sample_manager_inst.add_one_monitor(fifo_monitor_1082);
    sample_manager_inst.add_one_monitor(fifo_monitor_1083);
    sample_manager_inst.add_one_monitor(fifo_monitor_1084);
    sample_manager_inst.add_one_monitor(fifo_monitor_1085);
    sample_manager_inst.add_one_monitor(fifo_monitor_1086);
    sample_manager_inst.add_one_monitor(fifo_monitor_1087);
    sample_manager_inst.add_one_monitor(fifo_monitor_1088);
    sample_manager_inst.add_one_monitor(fifo_monitor_1089);
    sample_manager_inst.add_one_monitor(fifo_monitor_1090);
    sample_manager_inst.add_one_monitor(fifo_monitor_1091);
    sample_manager_inst.add_one_monitor(fifo_monitor_1092);
    sample_manager_inst.add_one_monitor(fifo_monitor_1093);
    sample_manager_inst.add_one_monitor(fifo_monitor_1094);
    sample_manager_inst.add_one_monitor(fifo_monitor_1095);
    sample_manager_inst.add_one_monitor(fifo_monitor_1096);
    sample_manager_inst.add_one_monitor(fifo_monitor_1097);
    sample_manager_inst.add_one_monitor(fifo_monitor_1098);
    sample_manager_inst.add_one_monitor(fifo_monitor_1099);
    sample_manager_inst.add_one_monitor(fifo_monitor_1100);
    sample_manager_inst.add_one_monitor(fifo_monitor_1101);
    sample_manager_inst.add_one_monitor(fifo_monitor_1102);
    sample_manager_inst.add_one_monitor(fifo_monitor_1103);
    sample_manager_inst.add_one_monitor(fifo_monitor_1104);
    sample_manager_inst.add_one_monitor(fifo_monitor_1105);
    sample_manager_inst.add_one_monitor(fifo_monitor_1106);
    sample_manager_inst.add_one_monitor(fifo_monitor_1107);
    sample_manager_inst.add_one_monitor(fifo_monitor_1108);
    sample_manager_inst.add_one_monitor(fifo_monitor_1109);
    sample_manager_inst.add_one_monitor(fifo_monitor_1110);
    sample_manager_inst.add_one_monitor(fifo_monitor_1111);
    sample_manager_inst.add_one_monitor(fifo_monitor_1112);
    sample_manager_inst.add_one_monitor(fifo_monitor_1113);
    sample_manager_inst.add_one_monitor(fifo_monitor_1114);
    sample_manager_inst.add_one_monitor(fifo_monitor_1115);
    sample_manager_inst.add_one_monitor(fifo_monitor_1116);
    sample_manager_inst.add_one_monitor(fifo_monitor_1117);
    sample_manager_inst.add_one_monitor(fifo_monitor_1118);
    sample_manager_inst.add_one_monitor(fifo_monitor_1119);
    sample_manager_inst.add_one_monitor(fifo_monitor_1120);
    sample_manager_inst.add_one_monitor(fifo_monitor_1121);
    sample_manager_inst.add_one_monitor(fifo_monitor_1122);
    sample_manager_inst.add_one_monitor(fifo_monitor_1123);
    sample_manager_inst.add_one_monitor(fifo_monitor_1124);
    sample_manager_inst.add_one_monitor(fifo_monitor_1125);
    sample_manager_inst.add_one_monitor(fifo_monitor_1126);
    sample_manager_inst.add_one_monitor(fifo_monitor_1127);
    sample_manager_inst.add_one_monitor(fifo_monitor_1128);
    sample_manager_inst.add_one_monitor(fifo_monitor_1129);
    sample_manager_inst.add_one_monitor(fifo_monitor_1130);
    sample_manager_inst.add_one_monitor(fifo_monitor_1131);
    sample_manager_inst.add_one_monitor(fifo_monitor_1132);
    sample_manager_inst.add_one_monitor(fifo_monitor_1133);
    sample_manager_inst.add_one_monitor(fifo_monitor_1134);
    sample_manager_inst.add_one_monitor(fifo_monitor_1135);
    sample_manager_inst.add_one_monitor(fifo_monitor_1136);
    sample_manager_inst.add_one_monitor(fifo_monitor_1137);
    sample_manager_inst.add_one_monitor(fifo_monitor_1138);
    sample_manager_inst.add_one_monitor(fifo_monitor_1139);
    sample_manager_inst.add_one_monitor(fifo_monitor_1140);
    sample_manager_inst.add_one_monitor(fifo_monitor_1141);
    sample_manager_inst.add_one_monitor(fifo_monitor_1142);
    sample_manager_inst.add_one_monitor(fifo_monitor_1143);
    sample_manager_inst.add_one_monitor(fifo_monitor_1144);
    sample_manager_inst.add_one_monitor(fifo_monitor_1145);
    sample_manager_inst.add_one_monitor(fifo_monitor_1146);
    sample_manager_inst.add_one_monitor(fifo_monitor_1147);
    sample_manager_inst.add_one_monitor(fifo_monitor_1148);
    sample_manager_inst.add_one_monitor(fifo_monitor_1149);
    sample_manager_inst.add_one_monitor(fifo_monitor_1150);
    sample_manager_inst.add_one_monitor(fifo_monitor_1151);
    sample_manager_inst.add_one_monitor(fifo_monitor_1152);
    sample_manager_inst.add_one_monitor(fifo_monitor_1153);
    sample_manager_inst.add_one_monitor(fifo_monitor_1154);
    sample_manager_inst.add_one_monitor(fifo_monitor_1155);
    sample_manager_inst.add_one_monitor(fifo_monitor_1156);
    sample_manager_inst.add_one_monitor(fifo_monitor_1157);
    sample_manager_inst.add_one_monitor(fifo_monitor_1158);
    sample_manager_inst.add_one_monitor(fifo_monitor_1159);
    sample_manager_inst.add_one_monitor(fifo_monitor_1160);
    sample_manager_inst.add_one_monitor(fifo_monitor_1161);
    sample_manager_inst.add_one_monitor(fifo_monitor_1162);
    sample_manager_inst.add_one_monitor(fifo_monitor_1163);
    sample_manager_inst.add_one_monitor(fifo_monitor_1164);
    sample_manager_inst.add_one_monitor(fifo_monitor_1165);
    sample_manager_inst.add_one_monitor(fifo_monitor_1166);
    sample_manager_inst.add_one_monitor(fifo_monitor_1167);
    sample_manager_inst.add_one_monitor(fifo_monitor_1168);
    sample_manager_inst.add_one_monitor(fifo_monitor_1169);
    sample_manager_inst.add_one_monitor(fifo_monitor_1170);
    sample_manager_inst.add_one_monitor(fifo_monitor_1171);
    sample_manager_inst.add_one_monitor(fifo_monitor_1172);
    sample_manager_inst.add_one_monitor(fifo_monitor_1173);
    sample_manager_inst.add_one_monitor(fifo_monitor_1174);
    sample_manager_inst.add_one_monitor(fifo_monitor_1175);
    sample_manager_inst.add_one_monitor(fifo_monitor_1176);
    sample_manager_inst.add_one_monitor(fifo_monitor_1177);
    sample_manager_inst.add_one_monitor(fifo_monitor_1178);
    sample_manager_inst.add_one_monitor(fifo_monitor_1179);
    sample_manager_inst.add_one_monitor(fifo_monitor_1180);
    sample_manager_inst.add_one_monitor(fifo_monitor_1181);
    sample_manager_inst.add_one_monitor(fifo_monitor_1182);
    sample_manager_inst.add_one_monitor(fifo_monitor_1183);
    sample_manager_inst.add_one_monitor(fifo_monitor_1184);
    sample_manager_inst.add_one_monitor(fifo_monitor_1185);
    sample_manager_inst.add_one_monitor(fifo_monitor_1186);
    sample_manager_inst.add_one_monitor(fifo_monitor_1187);
    sample_manager_inst.add_one_monitor(fifo_monitor_1188);
    sample_manager_inst.add_one_monitor(fifo_monitor_1189);
    sample_manager_inst.add_one_monitor(fifo_monitor_1190);
    sample_manager_inst.add_one_monitor(fifo_monitor_1191);
    sample_manager_inst.add_one_monitor(fifo_monitor_1192);
    sample_manager_inst.add_one_monitor(fifo_monitor_1193);
    sample_manager_inst.add_one_monitor(fifo_monitor_1194);
    sample_manager_inst.add_one_monitor(fifo_monitor_1195);
    sample_manager_inst.add_one_monitor(fifo_monitor_1196);
    sample_manager_inst.add_one_monitor(fifo_monitor_1197);
    sample_manager_inst.add_one_monitor(fifo_monitor_1198);
    sample_manager_inst.add_one_monitor(fifo_monitor_1199);
    sample_manager_inst.add_one_monitor(fifo_monitor_1200);
    sample_manager_inst.add_one_monitor(fifo_monitor_1201);
    sample_manager_inst.add_one_monitor(fifo_monitor_1202);
    sample_manager_inst.add_one_monitor(fifo_monitor_1203);
    sample_manager_inst.add_one_monitor(fifo_monitor_1204);
    sample_manager_inst.add_one_monitor(fifo_monitor_1205);
    sample_manager_inst.add_one_monitor(fifo_monitor_1206);
    sample_manager_inst.add_one_monitor(fifo_monitor_1207);
    sample_manager_inst.add_one_monitor(fifo_monitor_1208);
    sample_manager_inst.add_one_monitor(fifo_monitor_1209);
    sample_manager_inst.add_one_monitor(fifo_monitor_1210);
    sample_manager_inst.add_one_monitor(fifo_monitor_1211);
    sample_manager_inst.add_one_monitor(fifo_monitor_1212);
    sample_manager_inst.add_one_monitor(fifo_monitor_1213);
    sample_manager_inst.add_one_monitor(fifo_monitor_1214);
    sample_manager_inst.add_one_monitor(fifo_monitor_1215);
    sample_manager_inst.add_one_monitor(fifo_monitor_1216);
    sample_manager_inst.add_one_monitor(fifo_monitor_1217);
    sample_manager_inst.add_one_monitor(fifo_monitor_1218);
    sample_manager_inst.add_one_monitor(fifo_monitor_1219);
    sample_manager_inst.add_one_monitor(fifo_monitor_1220);
    sample_manager_inst.add_one_monitor(fifo_monitor_1221);
    sample_manager_inst.add_one_monitor(fifo_monitor_1222);
    sample_manager_inst.add_one_monitor(fifo_monitor_1223);
    sample_manager_inst.add_one_monitor(fifo_monitor_1224);
    sample_manager_inst.add_one_monitor(fifo_monitor_1225);
    sample_manager_inst.add_one_monitor(fifo_monitor_1226);
    sample_manager_inst.add_one_monitor(fifo_monitor_1227);
    sample_manager_inst.add_one_monitor(fifo_monitor_1228);
    sample_manager_inst.add_one_monitor(fifo_monitor_1229);
    sample_manager_inst.add_one_monitor(fifo_monitor_1230);
    sample_manager_inst.add_one_monitor(fifo_monitor_1231);
    sample_manager_inst.add_one_monitor(fifo_monitor_1232);
    sample_manager_inst.add_one_monitor(fifo_monitor_1233);
    sample_manager_inst.add_one_monitor(fifo_monitor_1234);
    sample_manager_inst.add_one_monitor(fifo_monitor_1235);
    sample_manager_inst.add_one_monitor(fifo_monitor_1236);
    sample_manager_inst.add_one_monitor(fifo_monitor_1237);
    sample_manager_inst.add_one_monitor(fifo_monitor_1238);
    sample_manager_inst.add_one_monitor(fifo_monitor_1239);
    sample_manager_inst.add_one_monitor(fifo_monitor_1240);
    sample_manager_inst.add_one_monitor(fifo_monitor_1241);
    sample_manager_inst.add_one_monitor(fifo_monitor_1242);
    sample_manager_inst.add_one_monitor(fifo_monitor_1243);
    sample_manager_inst.add_one_monitor(fifo_monitor_1244);
    sample_manager_inst.add_one_monitor(fifo_monitor_1245);
    sample_manager_inst.add_one_monitor(fifo_monitor_1246);
    sample_manager_inst.add_one_monitor(fifo_monitor_1247);
    sample_manager_inst.add_one_monitor(fifo_monitor_1248);
    sample_manager_inst.add_one_monitor(fifo_monitor_1249);
    sample_manager_inst.add_one_monitor(fifo_monitor_1250);
    sample_manager_inst.add_one_monitor(fifo_monitor_1251);
    sample_manager_inst.add_one_monitor(fifo_monitor_1252);
    sample_manager_inst.add_one_monitor(fifo_monitor_1253);
    sample_manager_inst.add_one_monitor(fifo_monitor_1254);
    sample_manager_inst.add_one_monitor(fifo_monitor_1255);
    sample_manager_inst.add_one_monitor(fifo_monitor_1256);
    sample_manager_inst.add_one_monitor(fifo_monitor_1257);
    sample_manager_inst.add_one_monitor(fifo_monitor_1258);
    sample_manager_inst.add_one_monitor(fifo_monitor_1259);
    sample_manager_inst.add_one_monitor(fifo_monitor_1260);
    sample_manager_inst.add_one_monitor(fifo_monitor_1261);
    sample_manager_inst.add_one_monitor(fifo_monitor_1262);
    sample_manager_inst.add_one_monitor(fifo_monitor_1263);
    sample_manager_inst.add_one_monitor(fifo_monitor_1264);
    sample_manager_inst.add_one_monitor(fifo_monitor_1265);
    sample_manager_inst.add_one_monitor(fifo_monitor_1266);
    sample_manager_inst.add_one_monitor(fifo_monitor_1267);
    sample_manager_inst.add_one_monitor(fifo_monitor_1268);
    sample_manager_inst.add_one_monitor(fifo_monitor_1269);
    sample_manager_inst.add_one_monitor(fifo_monitor_1270);
    sample_manager_inst.add_one_monitor(fifo_monitor_1271);
    sample_manager_inst.add_one_monitor(fifo_monitor_1272);
    sample_manager_inst.add_one_monitor(fifo_monitor_1273);
    sample_manager_inst.add_one_monitor(fifo_monitor_1274);
    sample_manager_inst.add_one_monitor(fifo_monitor_1275);
    sample_manager_inst.add_one_monitor(fifo_monitor_1276);
    sample_manager_inst.add_one_monitor(fifo_monitor_1277);
    sample_manager_inst.add_one_monitor(fifo_monitor_1278);
    sample_manager_inst.add_one_monitor(fifo_monitor_1279);
    sample_manager_inst.add_one_monitor(fifo_monitor_1280);
    sample_manager_inst.add_one_monitor(fifo_monitor_1281);
    sample_manager_inst.add_one_monitor(fifo_monitor_1282);
    sample_manager_inst.add_one_monitor(fifo_monitor_1283);
    sample_manager_inst.add_one_monitor(fifo_monitor_1284);
    sample_manager_inst.add_one_monitor(fifo_monitor_1285);
    sample_manager_inst.add_one_monitor(fifo_monitor_1286);
    sample_manager_inst.add_one_monitor(fifo_monitor_1287);
    sample_manager_inst.add_one_monitor(fifo_monitor_1288);
    sample_manager_inst.add_one_monitor(fifo_monitor_1289);
    sample_manager_inst.add_one_monitor(fifo_monitor_1290);
    sample_manager_inst.add_one_monitor(fifo_monitor_1291);
    sample_manager_inst.add_one_monitor(fifo_monitor_1292);
    sample_manager_inst.add_one_monitor(fifo_monitor_1293);
    sample_manager_inst.add_one_monitor(fifo_monitor_1294);
    sample_manager_inst.add_one_monitor(fifo_monitor_1295);
    sample_manager_inst.add_one_monitor(fifo_monitor_1296);
    sample_manager_inst.add_one_monitor(fifo_monitor_1297);
    sample_manager_inst.add_one_monitor(fifo_monitor_1298);
    sample_manager_inst.add_one_monitor(fifo_monitor_1299);
    sample_manager_inst.add_one_monitor(fifo_monitor_1300);
    sample_manager_inst.add_one_monitor(fifo_monitor_1301);
    sample_manager_inst.add_one_monitor(fifo_monitor_1302);
    sample_manager_inst.add_one_monitor(fifo_monitor_1303);
    sample_manager_inst.add_one_monitor(fifo_monitor_1304);
    sample_manager_inst.add_one_monitor(fifo_monitor_1305);
    sample_manager_inst.add_one_monitor(fifo_monitor_1306);
    sample_manager_inst.add_one_monitor(fifo_monitor_1307);
    sample_manager_inst.add_one_monitor(fifo_monitor_1308);
    sample_manager_inst.add_one_monitor(fifo_monitor_1309);
    sample_manager_inst.add_one_monitor(fifo_monitor_1310);
    sample_manager_inst.add_one_monitor(fifo_monitor_1311);
    sample_manager_inst.add_one_monitor(fifo_monitor_1312);
    sample_manager_inst.add_one_monitor(fifo_monitor_1313);
    sample_manager_inst.add_one_monitor(fifo_monitor_1314);
    sample_manager_inst.add_one_monitor(fifo_monitor_1315);
    sample_manager_inst.add_one_monitor(fifo_monitor_1316);
    sample_manager_inst.add_one_monitor(fifo_monitor_1317);
    sample_manager_inst.add_one_monitor(fifo_monitor_1318);
    sample_manager_inst.add_one_monitor(fifo_monitor_1319);
    sample_manager_inst.add_one_monitor(fifo_monitor_1320);
    sample_manager_inst.add_one_monitor(fifo_monitor_1321);
    sample_manager_inst.add_one_monitor(fifo_monitor_1322);
    sample_manager_inst.add_one_monitor(fifo_monitor_1323);
    sample_manager_inst.add_one_monitor(fifo_monitor_1324);
    sample_manager_inst.add_one_monitor(fifo_monitor_1325);
    sample_manager_inst.add_one_monitor(fifo_monitor_1326);
    sample_manager_inst.add_one_monitor(fifo_monitor_1327);
    sample_manager_inst.add_one_monitor(fifo_monitor_1328);
    sample_manager_inst.add_one_monitor(fifo_monitor_1329);
    sample_manager_inst.add_one_monitor(fifo_monitor_1330);
    sample_manager_inst.add_one_monitor(fifo_monitor_1331);
    sample_manager_inst.add_one_monitor(fifo_monitor_1332);
    sample_manager_inst.add_one_monitor(fifo_monitor_1333);
    sample_manager_inst.add_one_monitor(fifo_monitor_1334);
    sample_manager_inst.add_one_monitor(fifo_monitor_1335);
    sample_manager_inst.add_one_monitor(fifo_monitor_1336);
    sample_manager_inst.add_one_monitor(fifo_monitor_1337);
    sample_manager_inst.add_one_monitor(fifo_monitor_1338);
    sample_manager_inst.add_one_monitor(fifo_monitor_1339);
    sample_manager_inst.add_one_monitor(fifo_monitor_1340);
    sample_manager_inst.add_one_monitor(fifo_monitor_1341);
    sample_manager_inst.add_one_monitor(fifo_monitor_1342);
    sample_manager_inst.add_one_monitor(fifo_monitor_1343);
    sample_manager_inst.add_one_monitor(fifo_monitor_1344);
    sample_manager_inst.add_one_monitor(fifo_monitor_1345);
    sample_manager_inst.add_one_monitor(fifo_monitor_1346);
    sample_manager_inst.add_one_monitor(fifo_monitor_1347);
    sample_manager_inst.add_one_monitor(fifo_monitor_1348);
    sample_manager_inst.add_one_monitor(fifo_monitor_1349);
    sample_manager_inst.add_one_monitor(fifo_monitor_1350);
    sample_manager_inst.add_one_monitor(fifo_monitor_1351);
    sample_manager_inst.add_one_monitor(fifo_monitor_1352);
    sample_manager_inst.add_one_monitor(fifo_monitor_1353);
    sample_manager_inst.add_one_monitor(fifo_monitor_1354);
    sample_manager_inst.add_one_monitor(fifo_monitor_1355);
    sample_manager_inst.add_one_monitor(fifo_monitor_1356);
    sample_manager_inst.add_one_monitor(fifo_monitor_1357);
    sample_manager_inst.add_one_monitor(fifo_monitor_1358);
    sample_manager_inst.add_one_monitor(fifo_monitor_1359);
    sample_manager_inst.add_one_monitor(fifo_monitor_1360);
    sample_manager_inst.add_one_monitor(fifo_monitor_1361);
    sample_manager_inst.add_one_monitor(fifo_monitor_1362);
    sample_manager_inst.add_one_monitor(fifo_monitor_1363);
    sample_manager_inst.add_one_monitor(fifo_monitor_1364);
    sample_manager_inst.add_one_monitor(fifo_monitor_1365);
    sample_manager_inst.add_one_monitor(fifo_monitor_1366);
    sample_manager_inst.add_one_monitor(fifo_monitor_1367);
    sample_manager_inst.add_one_monitor(fifo_monitor_1368);
    sample_manager_inst.add_one_monitor(fifo_monitor_1369);
    sample_manager_inst.add_one_monitor(fifo_monitor_1370);
    sample_manager_inst.add_one_monitor(fifo_monitor_1371);
    sample_manager_inst.add_one_monitor(fifo_monitor_1372);
    sample_manager_inst.add_one_monitor(fifo_monitor_1373);
    sample_manager_inst.add_one_monitor(fifo_monitor_1374);
    sample_manager_inst.add_one_monitor(fifo_monitor_1375);
    sample_manager_inst.add_one_monitor(fifo_monitor_1376);
    sample_manager_inst.add_one_monitor(fifo_monitor_1377);
    sample_manager_inst.add_one_monitor(fifo_monitor_1378);
    sample_manager_inst.add_one_monitor(fifo_monitor_1379);
    sample_manager_inst.add_one_monitor(fifo_monitor_1380);
    sample_manager_inst.add_one_monitor(fifo_monitor_1381);
    sample_manager_inst.add_one_monitor(fifo_monitor_1382);
    sample_manager_inst.add_one_monitor(fifo_monitor_1383);
    sample_manager_inst.add_one_monitor(fifo_monitor_1384);
    sample_manager_inst.add_one_monitor(fifo_monitor_1385);
    sample_manager_inst.add_one_monitor(fifo_monitor_1386);
    sample_manager_inst.add_one_monitor(fifo_monitor_1387);
    sample_manager_inst.add_one_monitor(fifo_monitor_1388);
    sample_manager_inst.add_one_monitor(fifo_monitor_1389);
    sample_manager_inst.add_one_monitor(fifo_monitor_1390);
    sample_manager_inst.add_one_monitor(fifo_monitor_1391);
    sample_manager_inst.add_one_monitor(fifo_monitor_1392);
    sample_manager_inst.add_one_monitor(fifo_monitor_1393);
    sample_manager_inst.add_one_monitor(fifo_monitor_1394);
    sample_manager_inst.add_one_monitor(fifo_monitor_1395);
    sample_manager_inst.add_one_monitor(fifo_monitor_1396);
    sample_manager_inst.add_one_monitor(fifo_monitor_1397);
    sample_manager_inst.add_one_monitor(fifo_monitor_1398);
    sample_manager_inst.add_one_monitor(fifo_monitor_1399);
    sample_manager_inst.add_one_monitor(fifo_monitor_1400);
    sample_manager_inst.add_one_monitor(fifo_monitor_1401);
    sample_manager_inst.add_one_monitor(fifo_monitor_1402);
    sample_manager_inst.add_one_monitor(fifo_monitor_1403);
    sample_manager_inst.add_one_monitor(fifo_monitor_1404);
    sample_manager_inst.add_one_monitor(fifo_monitor_1405);
    sample_manager_inst.add_one_monitor(fifo_monitor_1406);
    sample_manager_inst.add_one_monitor(fifo_monitor_1407);
    sample_manager_inst.add_one_monitor(fifo_monitor_1408);
    sample_manager_inst.add_one_monitor(fifo_monitor_1409);
    sample_manager_inst.add_one_monitor(fifo_monitor_1410);
    sample_manager_inst.add_one_monitor(fifo_monitor_1411);
    sample_manager_inst.add_one_monitor(fifo_monitor_1412);
    sample_manager_inst.add_one_monitor(fifo_monitor_1413);
    sample_manager_inst.add_one_monitor(fifo_monitor_1414);
    sample_manager_inst.add_one_monitor(fifo_monitor_1415);
    sample_manager_inst.add_one_monitor(fifo_monitor_1416);
    sample_manager_inst.add_one_monitor(fifo_monitor_1417);
    sample_manager_inst.add_one_monitor(fifo_monitor_1418);
    sample_manager_inst.add_one_monitor(fifo_monitor_1419);
    sample_manager_inst.add_one_monitor(fifo_monitor_1420);
    sample_manager_inst.add_one_monitor(fifo_monitor_1421);
    sample_manager_inst.add_one_monitor(fifo_monitor_1422);
    sample_manager_inst.add_one_monitor(fifo_monitor_1423);
    sample_manager_inst.add_one_monitor(fifo_monitor_1424);
    sample_manager_inst.add_one_monitor(fifo_monitor_1425);
    sample_manager_inst.add_one_monitor(fifo_monitor_1426);
    sample_manager_inst.add_one_monitor(fifo_monitor_1427);
    sample_manager_inst.add_one_monitor(fifo_monitor_1428);
    sample_manager_inst.add_one_monitor(fifo_monitor_1429);
    sample_manager_inst.add_one_monitor(fifo_monitor_1430);
    sample_manager_inst.add_one_monitor(fifo_monitor_1431);
    sample_manager_inst.add_one_monitor(fifo_monitor_1432);
    sample_manager_inst.add_one_monitor(fifo_monitor_1433);
    sample_manager_inst.add_one_monitor(fifo_monitor_1434);
    sample_manager_inst.add_one_monitor(fifo_monitor_1435);
    sample_manager_inst.add_one_monitor(fifo_monitor_1436);
    sample_manager_inst.add_one_monitor(fifo_monitor_1437);
    sample_manager_inst.add_one_monitor(fifo_monitor_1438);
    sample_manager_inst.add_one_monitor(fifo_monitor_1439);
    sample_manager_inst.add_one_monitor(fifo_monitor_1440);
    sample_manager_inst.add_one_monitor(fifo_monitor_1441);
    sample_manager_inst.add_one_monitor(fifo_monitor_1442);
    sample_manager_inst.add_one_monitor(fifo_monitor_1443);
    sample_manager_inst.add_one_monitor(fifo_monitor_1444);
    sample_manager_inst.add_one_monitor(fifo_monitor_1445);
    sample_manager_inst.add_one_monitor(fifo_monitor_1446);
    sample_manager_inst.add_one_monitor(fifo_monitor_1447);
    sample_manager_inst.add_one_monitor(fifo_monitor_1448);
    sample_manager_inst.add_one_monitor(fifo_monitor_1449);
    sample_manager_inst.add_one_monitor(fifo_monitor_1450);
    sample_manager_inst.add_one_monitor(fifo_monitor_1451);
    sample_manager_inst.add_one_monitor(fifo_monitor_1452);
    sample_manager_inst.add_one_monitor(fifo_monitor_1453);
    sample_manager_inst.add_one_monitor(fifo_monitor_1454);
    sample_manager_inst.add_one_monitor(fifo_monitor_1455);
    sample_manager_inst.add_one_monitor(fifo_monitor_1456);
    sample_manager_inst.add_one_monitor(fifo_monitor_1457);
    sample_manager_inst.add_one_monitor(fifo_monitor_1458);
    sample_manager_inst.add_one_monitor(fifo_monitor_1459);
    sample_manager_inst.add_one_monitor(fifo_monitor_1460);
    sample_manager_inst.add_one_monitor(fifo_monitor_1461);
    sample_manager_inst.add_one_monitor(fifo_monitor_1462);
    sample_manager_inst.add_one_monitor(fifo_monitor_1463);
    sample_manager_inst.add_one_monitor(fifo_monitor_1464);
    sample_manager_inst.add_one_monitor(fifo_monitor_1465);
    sample_manager_inst.add_one_monitor(fifo_monitor_1466);
    sample_manager_inst.add_one_monitor(fifo_monitor_1467);
    sample_manager_inst.add_one_monitor(fifo_monitor_1468);
    sample_manager_inst.add_one_monitor(fifo_monitor_1469);
    sample_manager_inst.add_one_monitor(fifo_monitor_1470);
    sample_manager_inst.add_one_monitor(fifo_monitor_1471);
    sample_manager_inst.add_one_monitor(fifo_monitor_1472);
    sample_manager_inst.add_one_monitor(fifo_monitor_1473);
    sample_manager_inst.add_one_monitor(fifo_monitor_1474);
    sample_manager_inst.add_one_monitor(fifo_monitor_1475);
    sample_manager_inst.add_one_monitor(fifo_monitor_1476);
    sample_manager_inst.add_one_monitor(fifo_monitor_1477);
    sample_manager_inst.add_one_monitor(fifo_monitor_1478);
    sample_manager_inst.add_one_monitor(fifo_monitor_1479);
    sample_manager_inst.add_one_monitor(fifo_monitor_1480);
    sample_manager_inst.add_one_monitor(fifo_monitor_1481);
    sample_manager_inst.add_one_monitor(fifo_monitor_1482);
    sample_manager_inst.add_one_monitor(fifo_monitor_1483);
    sample_manager_inst.add_one_monitor(fifo_monitor_1484);
    sample_manager_inst.add_one_monitor(fifo_monitor_1485);
    sample_manager_inst.add_one_monitor(fifo_monitor_1486);
    sample_manager_inst.add_one_monitor(fifo_monitor_1487);
    sample_manager_inst.add_one_monitor(fifo_monitor_1488);
    sample_manager_inst.add_one_monitor(fifo_monitor_1489);
    sample_manager_inst.add_one_monitor(fifo_monitor_1490);
    sample_manager_inst.add_one_monitor(fifo_monitor_1491);
    sample_manager_inst.add_one_monitor(fifo_monitor_1492);
    sample_manager_inst.add_one_monitor(fifo_monitor_1493);
    sample_manager_inst.add_one_monitor(fifo_monitor_1494);
    sample_manager_inst.add_one_monitor(fifo_monitor_1495);
    sample_manager_inst.add_one_monitor(fifo_monitor_1496);
    sample_manager_inst.add_one_monitor(fifo_monitor_1497);
    sample_manager_inst.add_one_monitor(fifo_monitor_1498);
    sample_manager_inst.add_one_monitor(fifo_monitor_1499);
    sample_manager_inst.add_one_monitor(fifo_monitor_1500);
    sample_manager_inst.add_one_monitor(fifo_monitor_1501);
    sample_manager_inst.add_one_monitor(fifo_monitor_1502);
    sample_manager_inst.add_one_monitor(fifo_monitor_1503);
    sample_manager_inst.add_one_monitor(fifo_monitor_1504);
    sample_manager_inst.add_one_monitor(fifo_monitor_1505);
    sample_manager_inst.add_one_monitor(fifo_monitor_1506);
    sample_manager_inst.add_one_monitor(fifo_monitor_1507);
    sample_manager_inst.add_one_monitor(fifo_monitor_1508);
    sample_manager_inst.add_one_monitor(fifo_monitor_1509);
    sample_manager_inst.add_one_monitor(fifo_monitor_1510);
    sample_manager_inst.add_one_monitor(fifo_monitor_1511);
    sample_manager_inst.add_one_monitor(fifo_monitor_1512);
    sample_manager_inst.add_one_monitor(fifo_monitor_1513);
    sample_manager_inst.add_one_monitor(fifo_monitor_1514);
    sample_manager_inst.add_one_monitor(fifo_monitor_1515);
    sample_manager_inst.add_one_monitor(fifo_monitor_1516);
    sample_manager_inst.add_one_monitor(fifo_monitor_1517);
    sample_manager_inst.add_one_monitor(fifo_monitor_1518);
    sample_manager_inst.add_one_monitor(fifo_monitor_1519);
    sample_manager_inst.add_one_monitor(fifo_monitor_1520);
    sample_manager_inst.add_one_monitor(fifo_monitor_1521);
    sample_manager_inst.add_one_monitor(fifo_monitor_1522);
    sample_manager_inst.add_one_monitor(fifo_monitor_1523);
    sample_manager_inst.add_one_monitor(fifo_monitor_1524);
    sample_manager_inst.add_one_monitor(fifo_monitor_1525);
    sample_manager_inst.add_one_monitor(fifo_monitor_1526);
    sample_manager_inst.add_one_monitor(fifo_monitor_1527);
    sample_manager_inst.add_one_monitor(fifo_monitor_1528);
    sample_manager_inst.add_one_monitor(fifo_monitor_1529);
    sample_manager_inst.add_one_monitor(fifo_monitor_1530);
    sample_manager_inst.add_one_monitor(fifo_monitor_1531);
    sample_manager_inst.add_one_monitor(fifo_monitor_1532);
    sample_manager_inst.add_one_monitor(fifo_monitor_1533);
    sample_manager_inst.add_one_monitor(fifo_monitor_1534);
    sample_manager_inst.add_one_monitor(fifo_monitor_1535);
    sample_manager_inst.add_one_monitor(fifo_monitor_1536);
    sample_manager_inst.add_one_monitor(fifo_monitor_1537);
    sample_manager_inst.add_one_monitor(fifo_monitor_1538);
    sample_manager_inst.add_one_monitor(fifo_monitor_1539);
    sample_manager_inst.add_one_monitor(fifo_monitor_1540);
    sample_manager_inst.add_one_monitor(fifo_monitor_1541);
    sample_manager_inst.add_one_monitor(fifo_monitor_1542);
    sample_manager_inst.add_one_monitor(fifo_monitor_1543);
    sample_manager_inst.add_one_monitor(fifo_monitor_1544);
    sample_manager_inst.add_one_monitor(fifo_monitor_1545);
    sample_manager_inst.add_one_monitor(fifo_monitor_1546);
    sample_manager_inst.add_one_monitor(fifo_monitor_1547);
    sample_manager_inst.add_one_monitor(fifo_monitor_1548);
    sample_manager_inst.add_one_monitor(fifo_monitor_1549);
    sample_manager_inst.add_one_monitor(fifo_monitor_1550);
    sample_manager_inst.add_one_monitor(fifo_monitor_1551);
    sample_manager_inst.add_one_monitor(fifo_monitor_1552);
    sample_manager_inst.add_one_monitor(fifo_monitor_1553);
    sample_manager_inst.add_one_monitor(fifo_monitor_1554);
    sample_manager_inst.add_one_monitor(fifo_monitor_1555);
    sample_manager_inst.add_one_monitor(fifo_monitor_1556);
    sample_manager_inst.add_one_monitor(fifo_monitor_1557);
    sample_manager_inst.add_one_monitor(fifo_monitor_1558);
    sample_manager_inst.add_one_monitor(fifo_monitor_1559);
    sample_manager_inst.add_one_monitor(fifo_monitor_1560);
    sample_manager_inst.add_one_monitor(fifo_monitor_1561);
    sample_manager_inst.add_one_monitor(fifo_monitor_1562);
    sample_manager_inst.add_one_monitor(fifo_monitor_1563);
    sample_manager_inst.add_one_monitor(fifo_monitor_1564);
    sample_manager_inst.add_one_monitor(fifo_monitor_1565);
    sample_manager_inst.add_one_monitor(fifo_monitor_1566);
    sample_manager_inst.add_one_monitor(fifo_monitor_1567);
    sample_manager_inst.add_one_monitor(fifo_monitor_1568);
    sample_manager_inst.add_one_monitor(fifo_monitor_1569);
    sample_manager_inst.add_one_monitor(fifo_monitor_1570);
    sample_manager_inst.add_one_monitor(fifo_monitor_1571);
    sample_manager_inst.add_one_monitor(fifo_monitor_1572);
    sample_manager_inst.add_one_monitor(fifo_monitor_1573);
    sample_manager_inst.add_one_monitor(fifo_monitor_1574);
    sample_manager_inst.add_one_monitor(fifo_monitor_1575);
    sample_manager_inst.add_one_monitor(fifo_monitor_1576);
    sample_manager_inst.add_one_monitor(fifo_monitor_1577);
    sample_manager_inst.add_one_monitor(fifo_monitor_1578);
    sample_manager_inst.add_one_monitor(fifo_monitor_1579);
    sample_manager_inst.add_one_monitor(fifo_monitor_1580);
    sample_manager_inst.add_one_monitor(fifo_monitor_1581);
    sample_manager_inst.add_one_monitor(fifo_monitor_1582);
    sample_manager_inst.add_one_monitor(fifo_monitor_1583);
    sample_manager_inst.add_one_monitor(fifo_monitor_1584);
    sample_manager_inst.add_one_monitor(fifo_monitor_1585);
    sample_manager_inst.add_one_monitor(fifo_monitor_1586);
    sample_manager_inst.add_one_monitor(fifo_monitor_1587);
    sample_manager_inst.add_one_monitor(fifo_monitor_1588);
    sample_manager_inst.add_one_monitor(fifo_monitor_1589);
    sample_manager_inst.add_one_monitor(fifo_monitor_1590);
    sample_manager_inst.add_one_monitor(fifo_monitor_1591);
    sample_manager_inst.add_one_monitor(fifo_monitor_1592);
    sample_manager_inst.add_one_monitor(fifo_monitor_1593);
    sample_manager_inst.add_one_monitor(fifo_monitor_1594);
    sample_manager_inst.add_one_monitor(fifo_monitor_1595);
    sample_manager_inst.add_one_monitor(fifo_monitor_1596);
    sample_manager_inst.add_one_monitor(fifo_monitor_1597);
    sample_manager_inst.add_one_monitor(fifo_monitor_1598);
    sample_manager_inst.add_one_monitor(fifo_monitor_1599);
    sample_manager_inst.add_one_monitor(fifo_monitor_1600);
    sample_manager_inst.add_one_monitor(fifo_monitor_1601);
    sample_manager_inst.add_one_monitor(fifo_monitor_1602);
    sample_manager_inst.add_one_monitor(fifo_monitor_1603);
    sample_manager_inst.add_one_monitor(fifo_monitor_1604);
    sample_manager_inst.add_one_monitor(fifo_monitor_1605);
    sample_manager_inst.add_one_monitor(fifo_monitor_1606);
    sample_manager_inst.add_one_monitor(fifo_monitor_1607);
    sample_manager_inst.add_one_monitor(fifo_monitor_1608);
    sample_manager_inst.add_one_monitor(fifo_monitor_1609);
    sample_manager_inst.add_one_monitor(fifo_monitor_1610);
    sample_manager_inst.add_one_monitor(fifo_monitor_1611);
    sample_manager_inst.add_one_monitor(fifo_monitor_1612);
    sample_manager_inst.add_one_monitor(fifo_monitor_1613);
    sample_manager_inst.add_one_monitor(fifo_monitor_1614);
    sample_manager_inst.add_one_monitor(fifo_monitor_1615);
    sample_manager_inst.add_one_monitor(fifo_monitor_1616);
    sample_manager_inst.add_one_monitor(fifo_monitor_1617);
    sample_manager_inst.add_one_monitor(fifo_monitor_1618);
    sample_manager_inst.add_one_monitor(fifo_monitor_1619);
    sample_manager_inst.add_one_monitor(fifo_monitor_1620);
    sample_manager_inst.add_one_monitor(fifo_monitor_1621);
    sample_manager_inst.add_one_monitor(fifo_monitor_1622);
    sample_manager_inst.add_one_monitor(fifo_monitor_1623);
    sample_manager_inst.add_one_monitor(fifo_monitor_1624);
    sample_manager_inst.add_one_monitor(fifo_monitor_1625);
    sample_manager_inst.add_one_monitor(fifo_monitor_1626);
    sample_manager_inst.add_one_monitor(fifo_monitor_1627);
    sample_manager_inst.add_one_monitor(fifo_monitor_1628);
    sample_manager_inst.add_one_monitor(fifo_monitor_1629);
    sample_manager_inst.add_one_monitor(fifo_monitor_1630);
    sample_manager_inst.add_one_monitor(fifo_monitor_1631);
    sample_manager_inst.add_one_monitor(fifo_monitor_1632);
    sample_manager_inst.add_one_monitor(fifo_monitor_1633);
    sample_manager_inst.add_one_monitor(fifo_monitor_1634);
    sample_manager_inst.add_one_monitor(fifo_monitor_1635);
    sample_manager_inst.add_one_monitor(fifo_monitor_1636);
    sample_manager_inst.add_one_monitor(fifo_monitor_1637);
    sample_manager_inst.add_one_monitor(fifo_monitor_1638);
    sample_manager_inst.add_one_monitor(fifo_monitor_1639);
    sample_manager_inst.add_one_monitor(fifo_monitor_1640);
    sample_manager_inst.add_one_monitor(fifo_monitor_1641);
    sample_manager_inst.add_one_monitor(fifo_monitor_1642);
    sample_manager_inst.add_one_monitor(fifo_monitor_1643);
    sample_manager_inst.add_one_monitor(fifo_monitor_1644);
    sample_manager_inst.add_one_monitor(fifo_monitor_1645);
    sample_manager_inst.add_one_monitor(fifo_monitor_1646);
    sample_manager_inst.add_one_monitor(fifo_monitor_1647);
    sample_manager_inst.add_one_monitor(fifo_monitor_1648);
    sample_manager_inst.add_one_monitor(fifo_monitor_1649);
    sample_manager_inst.add_one_monitor(fifo_monitor_1650);
    sample_manager_inst.add_one_monitor(fifo_monitor_1651);
    sample_manager_inst.add_one_monitor(fifo_monitor_1652);
    sample_manager_inst.add_one_monitor(fifo_monitor_1653);
    sample_manager_inst.add_one_monitor(fifo_monitor_1654);
    sample_manager_inst.add_one_monitor(fifo_monitor_1655);
    sample_manager_inst.add_one_monitor(fifo_monitor_1656);
    sample_manager_inst.add_one_monitor(fifo_monitor_1657);
    sample_manager_inst.add_one_monitor(fifo_monitor_1658);
    sample_manager_inst.add_one_monitor(fifo_monitor_1659);
    sample_manager_inst.add_one_monitor(fifo_monitor_1660);
    sample_manager_inst.add_one_monitor(fifo_monitor_1661);
    sample_manager_inst.add_one_monitor(fifo_monitor_1662);
    sample_manager_inst.add_one_monitor(fifo_monitor_1663);
    sample_manager_inst.add_one_monitor(fifo_monitor_1664);
    sample_manager_inst.add_one_monitor(fifo_monitor_1665);
    sample_manager_inst.add_one_monitor(fifo_monitor_1666);
    sample_manager_inst.add_one_monitor(fifo_monitor_1667);
    sample_manager_inst.add_one_monitor(fifo_monitor_1668);
    sample_manager_inst.add_one_monitor(fifo_monitor_1669);
    sample_manager_inst.add_one_monitor(fifo_monitor_1670);
    sample_manager_inst.add_one_monitor(fifo_monitor_1671);
    sample_manager_inst.add_one_monitor(fifo_monitor_1672);
    sample_manager_inst.add_one_monitor(fifo_monitor_1673);
    sample_manager_inst.add_one_monitor(fifo_monitor_1674);
    sample_manager_inst.add_one_monitor(fifo_monitor_1675);
    sample_manager_inst.add_one_monitor(fifo_monitor_1676);
    sample_manager_inst.add_one_monitor(fifo_monitor_1677);
    sample_manager_inst.add_one_monitor(fifo_monitor_1678);
    sample_manager_inst.add_one_monitor(fifo_monitor_1679);
    sample_manager_inst.add_one_monitor(fifo_monitor_1680);
    sample_manager_inst.add_one_monitor(fifo_monitor_1681);
    sample_manager_inst.add_one_monitor(fifo_monitor_1682);
    sample_manager_inst.add_one_monitor(fifo_monitor_1683);
    sample_manager_inst.add_one_monitor(fifo_monitor_1684);
    sample_manager_inst.add_one_monitor(fifo_monitor_1685);
    sample_manager_inst.add_one_monitor(fifo_monitor_1686);
    sample_manager_inst.add_one_monitor(fifo_monitor_1687);
    sample_manager_inst.add_one_monitor(fifo_monitor_1688);
    sample_manager_inst.add_one_monitor(fifo_monitor_1689);
    sample_manager_inst.add_one_monitor(fifo_monitor_1690);
    sample_manager_inst.add_one_monitor(fifo_monitor_1691);
    sample_manager_inst.add_one_monitor(fifo_monitor_1692);
    sample_manager_inst.add_one_monitor(fifo_monitor_1693);
    sample_manager_inst.add_one_monitor(fifo_monitor_1694);
    sample_manager_inst.add_one_monitor(fifo_monitor_1695);
    sample_manager_inst.add_one_monitor(fifo_monitor_1696);
    sample_manager_inst.add_one_monitor(fifo_monitor_1697);
    sample_manager_inst.add_one_monitor(fifo_monitor_1698);
    sample_manager_inst.add_one_monitor(fifo_monitor_1699);
    sample_manager_inst.add_one_monitor(fifo_monitor_1700);
    sample_manager_inst.add_one_monitor(fifo_monitor_1701);
    sample_manager_inst.add_one_monitor(fifo_monitor_1702);
    sample_manager_inst.add_one_monitor(fifo_monitor_1703);
    sample_manager_inst.add_one_monitor(fifo_monitor_1704);
    sample_manager_inst.add_one_monitor(fifo_monitor_1705);
    sample_manager_inst.add_one_monitor(fifo_monitor_1706);
    sample_manager_inst.add_one_monitor(fifo_monitor_1707);
    sample_manager_inst.add_one_monitor(fifo_monitor_1708);
    sample_manager_inst.add_one_monitor(fifo_monitor_1709);
    sample_manager_inst.add_one_monitor(fifo_monitor_1710);
    sample_manager_inst.add_one_monitor(fifo_monitor_1711);
    sample_manager_inst.add_one_monitor(fifo_monitor_1712);
    sample_manager_inst.add_one_monitor(fifo_monitor_1713);
    sample_manager_inst.add_one_monitor(fifo_monitor_1714);
    sample_manager_inst.add_one_monitor(fifo_monitor_1715);
    sample_manager_inst.add_one_monitor(fifo_monitor_1716);
    sample_manager_inst.add_one_monitor(fifo_monitor_1717);
    sample_manager_inst.add_one_monitor(fifo_monitor_1718);
    sample_manager_inst.add_one_monitor(fifo_monitor_1719);
    sample_manager_inst.add_one_monitor(fifo_monitor_1720);
    sample_manager_inst.add_one_monitor(fifo_monitor_1721);
    sample_manager_inst.add_one_monitor(fifo_monitor_1722);
    sample_manager_inst.add_one_monitor(fifo_monitor_1723);
    sample_manager_inst.add_one_monitor(fifo_monitor_1724);
    sample_manager_inst.add_one_monitor(fifo_monitor_1725);
    sample_manager_inst.add_one_monitor(fifo_monitor_1726);
    sample_manager_inst.add_one_monitor(fifo_monitor_1727);
    sample_manager_inst.add_one_monitor(fifo_monitor_1728);
    sample_manager_inst.add_one_monitor(fifo_monitor_1729);
    sample_manager_inst.add_one_monitor(fifo_monitor_1730);
    sample_manager_inst.add_one_monitor(fifo_monitor_1731);
    sample_manager_inst.add_one_monitor(fifo_monitor_1732);
    sample_manager_inst.add_one_monitor(fifo_monitor_1733);
    sample_manager_inst.add_one_monitor(fifo_monitor_1734);
    sample_manager_inst.add_one_monitor(fifo_monitor_1735);
    sample_manager_inst.add_one_monitor(fifo_monitor_1736);
    sample_manager_inst.add_one_monitor(fifo_monitor_1737);
    sample_manager_inst.add_one_monitor(fifo_monitor_1738);
    sample_manager_inst.add_one_monitor(fifo_monitor_1739);
    sample_manager_inst.add_one_monitor(fifo_monitor_1740);
    sample_manager_inst.add_one_monitor(fifo_monitor_1741);
    sample_manager_inst.add_one_monitor(fifo_monitor_1742);
    sample_manager_inst.add_one_monitor(fifo_monitor_1743);
    sample_manager_inst.add_one_monitor(fifo_monitor_1744);
    sample_manager_inst.add_one_monitor(fifo_monitor_1745);
    sample_manager_inst.add_one_monitor(fifo_monitor_1746);
    sample_manager_inst.add_one_monitor(fifo_monitor_1747);
    sample_manager_inst.add_one_monitor(fifo_monitor_1748);
    sample_manager_inst.add_one_monitor(fifo_monitor_1749);
    sample_manager_inst.add_one_monitor(fifo_monitor_1750);
    sample_manager_inst.add_one_monitor(fifo_monitor_1751);
    sample_manager_inst.add_one_monitor(fifo_monitor_1752);
    sample_manager_inst.add_one_monitor(fifo_monitor_1753);
    sample_manager_inst.add_one_monitor(fifo_monitor_1754);
    sample_manager_inst.add_one_monitor(fifo_monitor_1755);
    sample_manager_inst.add_one_monitor(fifo_monitor_1756);
    sample_manager_inst.add_one_monitor(fifo_monitor_1757);
    sample_manager_inst.add_one_monitor(fifo_monitor_1758);
    sample_manager_inst.add_one_monitor(fifo_monitor_1759);
    sample_manager_inst.add_one_monitor(fifo_monitor_1760);
    sample_manager_inst.add_one_monitor(fifo_monitor_1761);
    sample_manager_inst.add_one_monitor(fifo_monitor_1762);
    sample_manager_inst.add_one_monitor(fifo_monitor_1763);
    sample_manager_inst.add_one_monitor(fifo_monitor_1764);
    sample_manager_inst.add_one_monitor(fifo_monitor_1765);
    sample_manager_inst.add_one_monitor(fifo_monitor_1766);
    sample_manager_inst.add_one_monitor(fifo_monitor_1767);
    sample_manager_inst.add_one_monitor(fifo_monitor_1768);
    sample_manager_inst.add_one_monitor(fifo_monitor_1769);
    sample_manager_inst.add_one_monitor(fifo_monitor_1770);
    sample_manager_inst.add_one_monitor(fifo_monitor_1771);
    sample_manager_inst.add_one_monitor(fifo_monitor_1772);
    sample_manager_inst.add_one_monitor(fifo_monitor_1773);
    sample_manager_inst.add_one_monitor(fifo_monitor_1774);
    sample_manager_inst.add_one_monitor(fifo_monitor_1775);
    sample_manager_inst.add_one_monitor(fifo_monitor_1776);
    sample_manager_inst.add_one_monitor(fifo_monitor_1777);
    sample_manager_inst.add_one_monitor(fifo_monitor_1778);
    sample_manager_inst.add_one_monitor(fifo_monitor_1779);
    sample_manager_inst.add_one_monitor(fifo_monitor_1780);
    sample_manager_inst.add_one_monitor(fifo_monitor_1781);
    sample_manager_inst.add_one_monitor(fifo_monitor_1782);
    sample_manager_inst.add_one_monitor(fifo_monitor_1783);
    sample_manager_inst.add_one_monitor(fifo_monitor_1784);
    sample_manager_inst.add_one_monitor(fifo_monitor_1785);
    sample_manager_inst.add_one_monitor(fifo_monitor_1786);
    sample_manager_inst.add_one_monitor(fifo_monitor_1787);
    sample_manager_inst.add_one_monitor(fifo_monitor_1788);
    sample_manager_inst.add_one_monitor(fifo_monitor_1789);
    sample_manager_inst.add_one_monitor(fifo_monitor_1790);
    sample_manager_inst.add_one_monitor(fifo_monitor_1791);
    sample_manager_inst.add_one_monitor(fifo_monitor_1792);
    sample_manager_inst.add_one_monitor(fifo_monitor_1793);
    sample_manager_inst.add_one_monitor(fifo_monitor_1794);
    sample_manager_inst.add_one_monitor(fifo_monitor_1795);
    sample_manager_inst.add_one_monitor(fifo_monitor_1796);
    sample_manager_inst.add_one_monitor(fifo_monitor_1797);
    sample_manager_inst.add_one_monitor(fifo_monitor_1798);
    sample_manager_inst.add_one_monitor(fifo_monitor_1799);
    sample_manager_inst.add_one_monitor(fifo_monitor_1800);
    sample_manager_inst.add_one_monitor(fifo_monitor_1801);
    sample_manager_inst.add_one_monitor(fifo_monitor_1802);
    sample_manager_inst.add_one_monitor(fifo_monitor_1803);
    sample_manager_inst.add_one_monitor(fifo_monitor_1804);
    sample_manager_inst.add_one_monitor(fifo_monitor_1805);
    sample_manager_inst.add_one_monitor(fifo_monitor_1806);
    sample_manager_inst.add_one_monitor(fifo_monitor_1807);
    sample_manager_inst.add_one_monitor(fifo_monitor_1808);
    sample_manager_inst.add_one_monitor(fifo_monitor_1809);
    sample_manager_inst.add_one_monitor(fifo_monitor_1810);
    sample_manager_inst.add_one_monitor(fifo_monitor_1811);
    sample_manager_inst.add_one_monitor(fifo_monitor_1812);
    sample_manager_inst.add_one_monitor(fifo_monitor_1813);
    sample_manager_inst.add_one_monitor(fifo_monitor_1814);
    sample_manager_inst.add_one_monitor(fifo_monitor_1815);
    sample_manager_inst.add_one_monitor(fifo_monitor_1816);
    sample_manager_inst.add_one_monitor(fifo_monitor_1817);
    sample_manager_inst.add_one_monitor(fifo_monitor_1818);
    sample_manager_inst.add_one_monitor(fifo_monitor_1819);
    sample_manager_inst.add_one_monitor(fifo_monitor_1820);
    sample_manager_inst.add_one_monitor(fifo_monitor_1821);
    sample_manager_inst.add_one_monitor(fifo_monitor_1822);
    sample_manager_inst.add_one_monitor(fifo_monitor_1823);
    sample_manager_inst.add_one_monitor(fifo_monitor_1824);
    sample_manager_inst.add_one_monitor(fifo_monitor_1825);
    sample_manager_inst.add_one_monitor(fifo_monitor_1826);
    sample_manager_inst.add_one_monitor(fifo_monitor_1827);
    sample_manager_inst.add_one_monitor(fifo_monitor_1828);
    sample_manager_inst.add_one_monitor(fifo_monitor_1829);
    sample_manager_inst.add_one_monitor(fifo_monitor_1830);
    sample_manager_inst.add_one_monitor(fifo_monitor_1831);
    sample_manager_inst.add_one_monitor(fifo_monitor_1832);
    sample_manager_inst.add_one_monitor(fifo_monitor_1833);
    sample_manager_inst.add_one_monitor(fifo_monitor_1834);
    sample_manager_inst.add_one_monitor(fifo_monitor_1835);
    sample_manager_inst.add_one_monitor(fifo_monitor_1836);
    sample_manager_inst.add_one_monitor(fifo_monitor_1837);
    sample_manager_inst.add_one_monitor(fifo_monitor_1838);
    sample_manager_inst.add_one_monitor(fifo_monitor_1839);
    sample_manager_inst.add_one_monitor(fifo_monitor_1840);
    sample_manager_inst.add_one_monitor(fifo_monitor_1841);
    sample_manager_inst.add_one_monitor(fifo_monitor_1842);
    sample_manager_inst.add_one_monitor(fifo_monitor_1843);
    sample_manager_inst.add_one_monitor(fifo_monitor_1844);
    sample_manager_inst.add_one_monitor(fifo_monitor_1845);
    sample_manager_inst.add_one_monitor(fifo_monitor_1846);
    sample_manager_inst.add_one_monitor(fifo_monitor_1847);
    sample_manager_inst.add_one_monitor(fifo_monitor_1848);
    sample_manager_inst.add_one_monitor(fifo_monitor_1849);
    sample_manager_inst.add_one_monitor(fifo_monitor_1850);
    sample_manager_inst.add_one_monitor(fifo_monitor_1851);
    sample_manager_inst.add_one_monitor(fifo_monitor_1852);
    sample_manager_inst.add_one_monitor(fifo_monitor_1853);
    sample_manager_inst.add_one_monitor(fifo_monitor_1854);
    sample_manager_inst.add_one_monitor(fifo_monitor_1855);
    sample_manager_inst.add_one_monitor(fifo_monitor_1856);
    sample_manager_inst.add_one_monitor(fifo_monitor_1857);
    sample_manager_inst.add_one_monitor(fifo_monitor_1858);
    sample_manager_inst.add_one_monitor(fifo_monitor_1859);
    sample_manager_inst.add_one_monitor(fifo_monitor_1860);
    sample_manager_inst.add_one_monitor(fifo_monitor_1861);
    sample_manager_inst.add_one_monitor(fifo_monitor_1862);
    sample_manager_inst.add_one_monitor(fifo_monitor_1863);
    sample_manager_inst.add_one_monitor(fifo_monitor_1864);
    sample_manager_inst.add_one_monitor(fifo_monitor_1865);
    sample_manager_inst.add_one_monitor(fifo_monitor_1866);
    sample_manager_inst.add_one_monitor(fifo_monitor_1867);
    sample_manager_inst.add_one_monitor(fifo_monitor_1868);
    sample_manager_inst.add_one_monitor(fifo_monitor_1869);
    sample_manager_inst.add_one_monitor(fifo_monitor_1870);
    sample_manager_inst.add_one_monitor(fifo_monitor_1871);
    sample_manager_inst.add_one_monitor(fifo_monitor_1872);
    sample_manager_inst.add_one_monitor(fifo_monitor_1873);
    sample_manager_inst.add_one_monitor(fifo_monitor_1874);
    sample_manager_inst.add_one_monitor(fifo_monitor_1875);
    sample_manager_inst.add_one_monitor(fifo_monitor_1876);
    sample_manager_inst.add_one_monitor(fifo_monitor_1877);
    sample_manager_inst.add_one_monitor(fifo_monitor_1878);
    sample_manager_inst.add_one_monitor(fifo_monitor_1879);
    sample_manager_inst.add_one_monitor(fifo_monitor_1880);
    sample_manager_inst.add_one_monitor(fifo_monitor_1881);
    sample_manager_inst.add_one_monitor(fifo_monitor_1882);
    sample_manager_inst.add_one_monitor(fifo_monitor_1883);
    sample_manager_inst.add_one_monitor(fifo_monitor_1884);
    sample_manager_inst.add_one_monitor(fifo_monitor_1885);
    sample_manager_inst.add_one_monitor(fifo_monitor_1886);
    sample_manager_inst.add_one_monitor(fifo_monitor_1887);
    sample_manager_inst.add_one_monitor(fifo_monitor_1888);
    sample_manager_inst.add_one_monitor(fifo_monitor_1889);
    sample_manager_inst.add_one_monitor(fifo_monitor_1890);
    sample_manager_inst.add_one_monitor(fifo_monitor_1891);
    sample_manager_inst.add_one_monitor(fifo_monitor_1892);
    sample_manager_inst.add_one_monitor(fifo_monitor_1893);
    sample_manager_inst.add_one_monitor(fifo_monitor_1894);
    sample_manager_inst.add_one_monitor(fifo_monitor_1895);
    sample_manager_inst.add_one_monitor(fifo_monitor_1896);
    sample_manager_inst.add_one_monitor(fifo_monitor_1897);
    sample_manager_inst.add_one_monitor(fifo_monitor_1898);
    sample_manager_inst.add_one_monitor(fifo_monitor_1899);
    sample_manager_inst.add_one_monitor(fifo_monitor_1900);
    sample_manager_inst.add_one_monitor(fifo_monitor_1901);
    sample_manager_inst.add_one_monitor(fifo_monitor_1902);
    sample_manager_inst.add_one_monitor(fifo_monitor_1903);
    sample_manager_inst.add_one_monitor(fifo_monitor_1904);
    sample_manager_inst.add_one_monitor(fifo_monitor_1905);
    sample_manager_inst.add_one_monitor(fifo_monitor_1906);
    sample_manager_inst.add_one_monitor(fifo_monitor_1907);
    sample_manager_inst.add_one_monitor(fifo_monitor_1908);
    sample_manager_inst.add_one_monitor(fifo_monitor_1909);
    sample_manager_inst.add_one_monitor(fifo_monitor_1910);
    sample_manager_inst.add_one_monitor(fifo_monitor_1911);
    sample_manager_inst.add_one_monitor(fifo_monitor_1912);
    sample_manager_inst.add_one_monitor(fifo_monitor_1913);
    sample_manager_inst.add_one_monitor(fifo_monitor_1914);
    sample_manager_inst.add_one_monitor(fifo_monitor_1915);
    sample_manager_inst.add_one_monitor(fifo_monitor_1916);
    sample_manager_inst.add_one_monitor(fifo_monitor_1917);
    sample_manager_inst.add_one_monitor(fifo_monitor_1918);
    sample_manager_inst.add_one_monitor(fifo_monitor_1919);
    sample_manager_inst.add_one_monitor(fifo_monitor_1920);
    sample_manager_inst.add_one_monitor(fifo_monitor_1921);
    sample_manager_inst.add_one_monitor(fifo_monitor_1922);
    sample_manager_inst.add_one_monitor(fifo_monitor_1923);
    sample_manager_inst.add_one_monitor(fifo_monitor_1924);
    sample_manager_inst.add_one_monitor(fifo_monitor_1925);
    sample_manager_inst.add_one_monitor(fifo_monitor_1926);
    sample_manager_inst.add_one_monitor(fifo_monitor_1927);
    sample_manager_inst.add_one_monitor(fifo_monitor_1928);
    sample_manager_inst.add_one_monitor(fifo_monitor_1929);
    sample_manager_inst.add_one_monitor(fifo_monitor_1930);
    sample_manager_inst.add_one_monitor(fifo_monitor_1931);
    sample_manager_inst.add_one_monitor(fifo_monitor_1932);
    sample_manager_inst.add_one_monitor(fifo_monitor_1933);
    sample_manager_inst.add_one_monitor(fifo_monitor_1934);
    sample_manager_inst.add_one_monitor(fifo_monitor_1935);
    sample_manager_inst.add_one_monitor(fifo_monitor_1936);
    sample_manager_inst.add_one_monitor(fifo_monitor_1937);
    sample_manager_inst.add_one_monitor(fifo_monitor_1938);
    sample_manager_inst.add_one_monitor(fifo_monitor_1939);
    sample_manager_inst.add_one_monitor(fifo_monitor_1940);
    sample_manager_inst.add_one_monitor(fifo_monitor_1941);
    sample_manager_inst.add_one_monitor(fifo_monitor_1942);
    sample_manager_inst.add_one_monitor(fifo_monitor_1943);
    sample_manager_inst.add_one_monitor(fifo_monitor_1944);
    sample_manager_inst.add_one_monitor(fifo_monitor_1945);
    sample_manager_inst.add_one_monitor(fifo_monitor_1946);
    sample_manager_inst.add_one_monitor(fifo_monitor_1947);
    sample_manager_inst.add_one_monitor(fifo_monitor_1948);
    sample_manager_inst.add_one_monitor(fifo_monitor_1949);
    sample_manager_inst.add_one_monitor(fifo_monitor_1950);
    sample_manager_inst.add_one_monitor(fifo_monitor_1951);
    sample_manager_inst.add_one_monitor(fifo_monitor_1952);
    sample_manager_inst.add_one_monitor(fifo_monitor_1953);
    sample_manager_inst.add_one_monitor(fifo_monitor_1954);
    sample_manager_inst.add_one_monitor(fifo_monitor_1955);
    sample_manager_inst.add_one_monitor(fifo_monitor_1956);
    sample_manager_inst.add_one_monitor(fifo_monitor_1957);
    sample_manager_inst.add_one_monitor(fifo_monitor_1958);
    sample_manager_inst.add_one_monitor(fifo_monitor_1959);
    sample_manager_inst.add_one_monitor(fifo_monitor_1960);
    sample_manager_inst.add_one_monitor(fifo_monitor_1961);
    sample_manager_inst.add_one_monitor(fifo_monitor_1962);
    sample_manager_inst.add_one_monitor(fifo_monitor_1963);
    sample_manager_inst.add_one_monitor(fifo_monitor_1964);
    sample_manager_inst.add_one_monitor(fifo_monitor_1965);
    sample_manager_inst.add_one_monitor(fifo_monitor_1966);
    sample_manager_inst.add_one_monitor(fifo_monitor_1967);
    sample_manager_inst.add_one_monitor(fifo_monitor_1968);
    sample_manager_inst.add_one_monitor(fifo_monitor_1969);
    sample_manager_inst.add_one_monitor(fifo_monitor_1970);
    sample_manager_inst.add_one_monitor(fifo_monitor_1971);
    sample_manager_inst.add_one_monitor(fifo_monitor_1972);
    sample_manager_inst.add_one_monitor(fifo_monitor_1973);
    sample_manager_inst.add_one_monitor(fifo_monitor_1974);
    sample_manager_inst.add_one_monitor(fifo_monitor_1975);
    sample_manager_inst.add_one_monitor(fifo_monitor_1976);
    sample_manager_inst.add_one_monitor(fifo_monitor_1977);
    sample_manager_inst.add_one_monitor(fifo_monitor_1978);
    sample_manager_inst.add_one_monitor(fifo_monitor_1979);
    sample_manager_inst.add_one_monitor(fifo_monitor_1980);
    sample_manager_inst.add_one_monitor(fifo_monitor_1981);
    sample_manager_inst.add_one_monitor(fifo_monitor_1982);
    sample_manager_inst.add_one_monitor(fifo_monitor_1983);
    sample_manager_inst.add_one_monitor(fifo_monitor_1984);
    sample_manager_inst.add_one_monitor(fifo_monitor_1985);
    sample_manager_inst.add_one_monitor(fifo_monitor_1986);
    sample_manager_inst.add_one_monitor(fifo_monitor_1987);
    sample_manager_inst.add_one_monitor(fifo_monitor_1988);
    sample_manager_inst.add_one_monitor(fifo_monitor_1989);
    sample_manager_inst.add_one_monitor(fifo_monitor_1990);
    sample_manager_inst.add_one_monitor(fifo_monitor_1991);
    sample_manager_inst.add_one_monitor(fifo_monitor_1992);
    sample_manager_inst.add_one_monitor(fifo_monitor_1993);
    sample_manager_inst.add_one_monitor(fifo_monitor_1994);
    sample_manager_inst.add_one_monitor(fifo_monitor_1995);
    sample_manager_inst.add_one_monitor(fifo_monitor_1996);
    sample_manager_inst.add_one_monitor(fifo_monitor_1997);
    sample_manager_inst.add_one_monitor(fifo_monitor_1998);
    sample_manager_inst.add_one_monitor(fifo_monitor_1999);
    sample_manager_inst.add_one_monitor(fifo_monitor_2000);
    sample_manager_inst.add_one_monitor(fifo_monitor_2001);
    sample_manager_inst.add_one_monitor(fifo_monitor_2002);
    sample_manager_inst.add_one_monitor(fifo_monitor_2003);
    sample_manager_inst.add_one_monitor(fifo_monitor_2004);
    sample_manager_inst.add_one_monitor(fifo_monitor_2005);
    sample_manager_inst.add_one_monitor(fifo_monitor_2006);
    sample_manager_inst.add_one_monitor(fifo_monitor_2007);
    sample_manager_inst.add_one_monitor(fifo_monitor_2008);
    sample_manager_inst.add_one_monitor(fifo_monitor_2009);
    sample_manager_inst.add_one_monitor(fifo_monitor_2010);
    sample_manager_inst.add_one_monitor(fifo_monitor_2011);
    sample_manager_inst.add_one_monitor(fifo_monitor_2012);
    sample_manager_inst.add_one_monitor(fifo_monitor_2013);
    sample_manager_inst.add_one_monitor(fifo_monitor_2014);
    sample_manager_inst.add_one_monitor(fifo_monitor_2015);
    sample_manager_inst.add_one_monitor(fifo_monitor_2016);
    sample_manager_inst.add_one_monitor(fifo_monitor_2017);
    sample_manager_inst.add_one_monitor(fifo_monitor_2018);
    sample_manager_inst.add_one_monitor(fifo_monitor_2019);
    sample_manager_inst.add_one_monitor(fifo_monitor_2020);
    sample_manager_inst.add_one_monitor(fifo_monitor_2021);
    sample_manager_inst.add_one_monitor(fifo_monitor_2022);
    sample_manager_inst.add_one_monitor(fifo_monitor_2023);
    sample_manager_inst.add_one_monitor(fifo_monitor_2024);
    sample_manager_inst.add_one_monitor(fifo_monitor_2025);
    sample_manager_inst.add_one_monitor(fifo_monitor_2026);
    sample_manager_inst.add_one_monitor(fifo_monitor_2027);
    sample_manager_inst.add_one_monitor(fifo_monitor_2028);
    sample_manager_inst.add_one_monitor(fifo_monitor_2029);
    sample_manager_inst.add_one_monitor(fifo_monitor_2030);
    sample_manager_inst.add_one_monitor(fifo_monitor_2031);
    sample_manager_inst.add_one_monitor(fifo_monitor_2032);
    sample_manager_inst.add_one_monitor(fifo_monitor_2033);
    sample_manager_inst.add_one_monitor(fifo_monitor_2034);
    sample_manager_inst.add_one_monitor(fifo_monitor_2035);
    sample_manager_inst.add_one_monitor(fifo_monitor_2036);
    sample_manager_inst.add_one_monitor(fifo_monitor_2037);
    sample_manager_inst.add_one_monitor(fifo_monitor_2038);
    sample_manager_inst.add_one_monitor(fifo_monitor_2039);
    sample_manager_inst.add_one_monitor(fifo_monitor_2040);
    sample_manager_inst.add_one_monitor(fifo_monitor_2041);
    sample_manager_inst.add_one_monitor(fifo_monitor_2042);
    sample_manager_inst.add_one_monitor(fifo_monitor_2043);
    sample_manager_inst.add_one_monitor(fifo_monitor_2044);
    sample_manager_inst.add_one_monitor(fifo_monitor_2045);
    sample_manager_inst.add_one_monitor(fifo_monitor_2046);
    sample_manager_inst.add_one_monitor(fifo_monitor_2047);
    sample_manager_inst.add_one_monitor(fifo_monitor_2048);
    sample_manager_inst.add_one_monitor(fifo_monitor_2049);
    sample_manager_inst.add_one_monitor(fifo_monitor_2050);
    sample_manager_inst.add_one_monitor(fifo_monitor_2051);
    sample_manager_inst.add_one_monitor(fifo_monitor_2052);
    sample_manager_inst.add_one_monitor(fifo_monitor_2053);
    sample_manager_inst.add_one_monitor(fifo_monitor_2054);
    sample_manager_inst.add_one_monitor(fifo_monitor_2055);
    sample_manager_inst.add_one_monitor(fifo_monitor_2056);
    sample_manager_inst.add_one_monitor(fifo_monitor_2057);
    sample_manager_inst.add_one_monitor(fifo_monitor_2058);
    sample_manager_inst.add_one_monitor(fifo_monitor_2059);
    sample_manager_inst.add_one_monitor(fifo_monitor_2060);
    sample_manager_inst.add_one_monitor(fifo_monitor_2061);
    sample_manager_inst.add_one_monitor(fifo_monitor_2062);
    sample_manager_inst.add_one_monitor(fifo_monitor_2063);
    sample_manager_inst.add_one_monitor(fifo_monitor_2064);
    sample_manager_inst.add_one_monitor(fifo_monitor_2065);
    sample_manager_inst.add_one_monitor(fifo_monitor_2066);
    sample_manager_inst.add_one_monitor(fifo_monitor_2067);
    sample_manager_inst.add_one_monitor(fifo_monitor_2068);
    sample_manager_inst.add_one_monitor(fifo_monitor_2069);
    sample_manager_inst.add_one_monitor(fifo_monitor_2070);
    sample_manager_inst.add_one_monitor(fifo_monitor_2071);
    sample_manager_inst.add_one_monitor(fifo_monitor_2072);
    sample_manager_inst.add_one_monitor(fifo_monitor_2073);
    sample_manager_inst.add_one_monitor(fifo_monitor_2074);
    sample_manager_inst.add_one_monitor(fifo_monitor_2075);
    sample_manager_inst.add_one_monitor(fifo_monitor_2076);
    sample_manager_inst.add_one_monitor(fifo_monitor_2077);
    sample_manager_inst.add_one_monitor(fifo_monitor_2078);
    sample_manager_inst.add_one_monitor(fifo_monitor_2079);
    sample_manager_inst.add_one_monitor(fifo_monitor_2080);
    sample_manager_inst.add_one_monitor(fifo_monitor_2081);
    sample_manager_inst.add_one_monitor(fifo_monitor_2082);
    sample_manager_inst.add_one_monitor(fifo_monitor_2083);
    sample_manager_inst.add_one_monitor(fifo_monitor_2084);
    sample_manager_inst.add_one_monitor(fifo_monitor_2085);
    sample_manager_inst.add_one_monitor(fifo_monitor_2086);
    sample_manager_inst.add_one_monitor(fifo_monitor_2087);
    sample_manager_inst.add_one_monitor(fifo_monitor_2088);
    sample_manager_inst.add_one_monitor(fifo_monitor_2089);
    sample_manager_inst.add_one_monitor(fifo_monitor_2090);
    sample_manager_inst.add_one_monitor(fifo_monitor_2091);
    sample_manager_inst.add_one_monitor(fifo_monitor_2092);
    sample_manager_inst.add_one_monitor(fifo_monitor_2093);
    sample_manager_inst.add_one_monitor(fifo_monitor_2094);
    sample_manager_inst.add_one_monitor(fifo_monitor_2095);
    sample_manager_inst.add_one_monitor(fifo_monitor_2096);
    sample_manager_inst.add_one_monitor(fifo_monitor_2097);
    sample_manager_inst.add_one_monitor(fifo_monitor_2098);
    sample_manager_inst.add_one_monitor(fifo_monitor_2099);
    sample_manager_inst.add_one_monitor(fifo_monitor_2100);
    sample_manager_inst.add_one_monitor(fifo_monitor_2101);
    sample_manager_inst.add_one_monitor(fifo_monitor_2102);
    sample_manager_inst.add_one_monitor(fifo_monitor_2103);
    sample_manager_inst.add_one_monitor(fifo_monitor_2104);
    sample_manager_inst.add_one_monitor(fifo_monitor_2105);
    sample_manager_inst.add_one_monitor(fifo_monitor_2106);
    sample_manager_inst.add_one_monitor(fifo_monitor_2107);
    sample_manager_inst.add_one_monitor(fifo_monitor_2108);
    sample_manager_inst.add_one_monitor(fifo_monitor_2109);
    sample_manager_inst.add_one_monitor(fifo_monitor_2110);
    sample_manager_inst.add_one_monitor(fifo_monitor_2111);
    sample_manager_inst.add_one_monitor(fifo_monitor_2112);
    sample_manager_inst.add_one_monitor(fifo_monitor_2113);
    sample_manager_inst.add_one_monitor(fifo_monitor_2114);
    sample_manager_inst.add_one_monitor(fifo_monitor_2115);
    sample_manager_inst.add_one_monitor(fifo_monitor_2116);
    sample_manager_inst.add_one_monitor(fifo_monitor_2117);
    sample_manager_inst.add_one_monitor(fifo_monitor_2118);
    sample_manager_inst.add_one_monitor(fifo_monitor_2119);
    sample_manager_inst.add_one_monitor(fifo_monitor_2120);
    sample_manager_inst.add_one_monitor(fifo_monitor_2121);
    sample_manager_inst.add_one_monitor(fifo_monitor_2122);
    sample_manager_inst.add_one_monitor(fifo_monitor_2123);
    sample_manager_inst.add_one_monitor(fifo_monitor_2124);
    sample_manager_inst.add_one_monitor(fifo_monitor_2125);
    sample_manager_inst.add_one_monitor(fifo_monitor_2126);
    sample_manager_inst.add_one_monitor(fifo_monitor_2127);
    sample_manager_inst.add_one_monitor(fifo_monitor_2128);
    sample_manager_inst.add_one_monitor(fifo_monitor_2129);
    sample_manager_inst.add_one_monitor(fifo_monitor_2130);
    sample_manager_inst.add_one_monitor(fifo_monitor_2131);
    sample_manager_inst.add_one_monitor(fifo_monitor_2132);
    sample_manager_inst.add_one_monitor(fifo_monitor_2133);
    sample_manager_inst.add_one_monitor(fifo_monitor_2134);
    sample_manager_inst.add_one_monitor(fifo_monitor_2135);
    sample_manager_inst.add_one_monitor(fifo_monitor_2136);
    sample_manager_inst.add_one_monitor(fifo_monitor_2137);
    sample_manager_inst.add_one_monitor(fifo_monitor_2138);
    sample_manager_inst.add_one_monitor(fifo_monitor_2139);
    sample_manager_inst.add_one_monitor(fifo_monitor_2140);
    sample_manager_inst.add_one_monitor(fifo_monitor_2141);
    sample_manager_inst.add_one_monitor(fifo_monitor_2142);
    sample_manager_inst.add_one_monitor(fifo_monitor_2143);
    sample_manager_inst.add_one_monitor(fifo_monitor_2144);
    sample_manager_inst.add_one_monitor(fifo_monitor_2145);
    sample_manager_inst.add_one_monitor(fifo_monitor_2146);
    sample_manager_inst.add_one_monitor(fifo_monitor_2147);
    sample_manager_inst.add_one_monitor(fifo_monitor_2148);
    sample_manager_inst.add_one_monitor(fifo_monitor_2149);
    sample_manager_inst.add_one_monitor(fifo_monitor_2150);
    sample_manager_inst.add_one_monitor(fifo_monitor_2151);
    sample_manager_inst.add_one_monitor(fifo_monitor_2152);
    sample_manager_inst.add_one_monitor(fifo_monitor_2153);
    sample_manager_inst.add_one_monitor(fifo_monitor_2154);
    sample_manager_inst.add_one_monitor(fifo_monitor_2155);
    sample_manager_inst.add_one_monitor(fifo_monitor_2156);
    sample_manager_inst.add_one_monitor(fifo_monitor_2157);
    sample_manager_inst.add_one_monitor(fifo_monitor_2158);
    sample_manager_inst.add_one_monitor(fifo_monitor_2159);
    sample_manager_inst.add_one_monitor(fifo_monitor_2160);
    sample_manager_inst.add_one_monitor(fifo_monitor_2161);
    sample_manager_inst.add_one_monitor(fifo_monitor_2162);
    sample_manager_inst.add_one_monitor(fifo_monitor_2163);
    sample_manager_inst.add_one_monitor(fifo_monitor_2164);
    sample_manager_inst.add_one_monitor(fifo_monitor_2165);
    sample_manager_inst.add_one_monitor(fifo_monitor_2166);
    sample_manager_inst.add_one_monitor(fifo_monitor_2167);
    sample_manager_inst.add_one_monitor(fifo_monitor_2168);
    sample_manager_inst.add_one_monitor(fifo_monitor_2169);
    sample_manager_inst.add_one_monitor(fifo_monitor_2170);
    sample_manager_inst.add_one_monitor(fifo_monitor_2171);
    sample_manager_inst.add_one_monitor(fifo_monitor_2172);
    sample_manager_inst.add_one_monitor(fifo_monitor_2173);
    sample_manager_inst.add_one_monitor(fifo_monitor_2174);
    sample_manager_inst.add_one_monitor(fifo_monitor_2175);
    sample_manager_inst.add_one_monitor(fifo_monitor_2176);
    sample_manager_inst.add_one_monitor(fifo_monitor_2177);
    sample_manager_inst.add_one_monitor(fifo_monitor_2178);
    sample_manager_inst.add_one_monitor(fifo_monitor_2179);
    sample_manager_inst.add_one_monitor(fifo_monitor_2180);
    sample_manager_inst.add_one_monitor(fifo_monitor_2181);
    sample_manager_inst.add_one_monitor(fifo_monitor_2182);
    sample_manager_inst.add_one_monitor(fifo_monitor_2183);
    sample_manager_inst.add_one_monitor(fifo_monitor_2184);
    sample_manager_inst.add_one_monitor(fifo_monitor_2185);
    sample_manager_inst.add_one_monitor(fifo_monitor_2186);
    sample_manager_inst.add_one_monitor(fifo_monitor_2187);
    sample_manager_inst.add_one_monitor(fifo_monitor_2188);
    sample_manager_inst.add_one_monitor(fifo_monitor_2189);
    sample_manager_inst.add_one_monitor(fifo_monitor_2190);
    sample_manager_inst.add_one_monitor(fifo_monitor_2191);
    sample_manager_inst.add_one_monitor(fifo_monitor_2192);
    sample_manager_inst.add_one_monitor(fifo_monitor_2193);
    sample_manager_inst.add_one_monitor(fifo_monitor_2194);
    sample_manager_inst.add_one_monitor(fifo_monitor_2195);
    sample_manager_inst.add_one_monitor(fifo_monitor_2196);
    sample_manager_inst.add_one_monitor(fifo_monitor_2197);
    sample_manager_inst.add_one_monitor(fifo_monitor_2198);
    sample_manager_inst.add_one_monitor(fifo_monitor_2199);
    sample_manager_inst.add_one_monitor(fifo_monitor_2200);
    sample_manager_inst.add_one_monitor(fifo_monitor_2201);
    sample_manager_inst.add_one_monitor(fifo_monitor_2202);
    sample_manager_inst.add_one_monitor(fifo_monitor_2203);
    sample_manager_inst.add_one_monitor(fifo_monitor_2204);
    sample_manager_inst.add_one_monitor(fifo_monitor_2205);
    sample_manager_inst.add_one_monitor(fifo_monitor_2206);
    sample_manager_inst.add_one_monitor(fifo_monitor_2207);
    sample_manager_inst.add_one_monitor(fifo_monitor_2208);
    sample_manager_inst.add_one_monitor(fifo_monitor_2209);
    sample_manager_inst.add_one_monitor(fifo_monitor_2210);
    sample_manager_inst.add_one_monitor(fifo_monitor_2211);
    sample_manager_inst.add_one_monitor(fifo_monitor_2212);
    sample_manager_inst.add_one_monitor(fifo_monitor_2213);
    sample_manager_inst.add_one_monitor(fifo_monitor_2214);
    sample_manager_inst.add_one_monitor(fifo_monitor_2215);
    sample_manager_inst.add_one_monitor(fifo_monitor_2216);
    sample_manager_inst.add_one_monitor(fifo_monitor_2217);
    sample_manager_inst.add_one_monitor(fifo_monitor_2218);
    sample_manager_inst.add_one_monitor(fifo_monitor_2219);
    sample_manager_inst.add_one_monitor(fifo_monitor_2220);
    sample_manager_inst.add_one_monitor(fifo_monitor_2221);
    sample_manager_inst.add_one_monitor(fifo_monitor_2222);
    sample_manager_inst.add_one_monitor(fifo_monitor_2223);
    sample_manager_inst.add_one_monitor(fifo_monitor_2224);
    sample_manager_inst.add_one_monitor(fifo_monitor_2225);
    sample_manager_inst.add_one_monitor(fifo_monitor_2226);
    sample_manager_inst.add_one_monitor(fifo_monitor_2227);
    sample_manager_inst.add_one_monitor(fifo_monitor_2228);
    sample_manager_inst.add_one_monitor(fifo_monitor_2229);
    sample_manager_inst.add_one_monitor(fifo_monitor_2230);
    sample_manager_inst.add_one_monitor(fifo_monitor_2231);
    sample_manager_inst.add_one_monitor(fifo_monitor_2232);
    sample_manager_inst.add_one_monitor(fifo_monitor_2233);
    sample_manager_inst.add_one_monitor(fifo_monitor_2234);
    sample_manager_inst.add_one_monitor(fifo_monitor_2235);
    sample_manager_inst.add_one_monitor(fifo_monitor_2236);
    sample_manager_inst.add_one_monitor(fifo_monitor_2237);
    sample_manager_inst.add_one_monitor(fifo_monitor_2238);
    sample_manager_inst.add_one_monitor(fifo_monitor_2239);
    sample_manager_inst.add_one_monitor(fifo_monitor_2240);
    sample_manager_inst.add_one_monitor(fifo_monitor_2241);
    sample_manager_inst.add_one_monitor(fifo_monitor_2242);
    sample_manager_inst.add_one_monitor(fifo_monitor_2243);
    sample_manager_inst.add_one_monitor(fifo_monitor_2244);
    sample_manager_inst.add_one_monitor(fifo_monitor_2245);
    sample_manager_inst.add_one_monitor(fifo_monitor_2246);
    sample_manager_inst.add_one_monitor(fifo_monitor_2247);
    sample_manager_inst.add_one_monitor(fifo_monitor_2248);
    sample_manager_inst.add_one_monitor(fifo_monitor_2249);
    sample_manager_inst.add_one_monitor(fifo_monitor_2250);
    sample_manager_inst.add_one_monitor(fifo_monitor_2251);
    sample_manager_inst.add_one_monitor(fifo_monitor_2252);
    sample_manager_inst.add_one_monitor(fifo_monitor_2253);
    sample_manager_inst.add_one_monitor(fifo_monitor_2254);
    sample_manager_inst.add_one_monitor(fifo_monitor_2255);
    sample_manager_inst.add_one_monitor(fifo_monitor_2256);
    sample_manager_inst.add_one_monitor(fifo_monitor_2257);
    sample_manager_inst.add_one_monitor(fifo_monitor_2258);
    sample_manager_inst.add_one_monitor(fifo_monitor_2259);
    sample_manager_inst.add_one_monitor(fifo_monitor_2260);
    sample_manager_inst.add_one_monitor(fifo_monitor_2261);
    sample_manager_inst.add_one_monitor(fifo_monitor_2262);
    sample_manager_inst.add_one_monitor(fifo_monitor_2263);
    sample_manager_inst.add_one_monitor(fifo_monitor_2264);
    sample_manager_inst.add_one_monitor(fifo_monitor_2265);
    sample_manager_inst.add_one_monitor(fifo_monitor_2266);
    sample_manager_inst.add_one_monitor(fifo_monitor_2267);
    sample_manager_inst.add_one_monitor(fifo_monitor_2268);
    sample_manager_inst.add_one_monitor(fifo_monitor_2269);
    sample_manager_inst.add_one_monitor(fifo_monitor_2270);
    sample_manager_inst.add_one_monitor(fifo_monitor_2271);
    sample_manager_inst.add_one_monitor(fifo_monitor_2272);
    sample_manager_inst.add_one_monitor(fifo_monitor_2273);
    sample_manager_inst.add_one_monitor(fifo_monitor_2274);
    sample_manager_inst.add_one_monitor(fifo_monitor_2275);
    sample_manager_inst.add_one_monitor(fifo_monitor_2276);
    sample_manager_inst.add_one_monitor(fifo_monitor_2277);
    sample_manager_inst.add_one_monitor(fifo_monitor_2278);
    sample_manager_inst.add_one_monitor(fifo_monitor_2279);
    sample_manager_inst.add_one_monitor(fifo_monitor_2280);
    sample_manager_inst.add_one_monitor(fifo_monitor_2281);
    sample_manager_inst.add_one_monitor(fifo_monitor_2282);
    sample_manager_inst.add_one_monitor(fifo_monitor_2283);
    sample_manager_inst.add_one_monitor(fifo_monitor_2284);
    sample_manager_inst.add_one_monitor(fifo_monitor_2285);
    sample_manager_inst.add_one_monitor(fifo_monitor_2286);
    sample_manager_inst.add_one_monitor(fifo_monitor_2287);
    sample_manager_inst.add_one_monitor(fifo_monitor_2288);
    sample_manager_inst.add_one_monitor(fifo_monitor_2289);
    sample_manager_inst.add_one_monitor(fifo_monitor_2290);
    sample_manager_inst.add_one_monitor(fifo_monitor_2291);
    sample_manager_inst.add_one_monitor(fifo_monitor_2292);
    sample_manager_inst.add_one_monitor(fifo_monitor_2293);
    sample_manager_inst.add_one_monitor(fifo_monitor_2294);
    sample_manager_inst.add_one_monitor(fifo_monitor_2295);
    sample_manager_inst.add_one_monitor(fifo_monitor_2296);
    sample_manager_inst.add_one_monitor(fifo_monitor_2297);
    sample_manager_inst.add_one_monitor(fifo_monitor_2298);
    sample_manager_inst.add_one_monitor(fifo_monitor_2299);
    sample_manager_inst.add_one_monitor(fifo_monitor_2300);
    sample_manager_inst.add_one_monitor(fifo_monitor_2301);
    sample_manager_inst.add_one_monitor(fifo_monitor_2302);
    sample_manager_inst.add_one_monitor(fifo_monitor_2303);
    sample_manager_inst.add_one_monitor(fifo_monitor_2304);
    sample_manager_inst.add_one_monitor(fifo_monitor_2305);
    sample_manager_inst.add_one_monitor(fifo_monitor_2306);
    sample_manager_inst.add_one_monitor(fifo_monitor_2307);
    sample_manager_inst.add_one_monitor(fifo_monitor_2308);
    sample_manager_inst.add_one_monitor(fifo_monitor_2309);
    sample_manager_inst.add_one_monitor(fifo_monitor_2310);
    sample_manager_inst.add_one_monitor(fifo_monitor_2311);
    sample_manager_inst.add_one_monitor(fifo_monitor_2312);
    sample_manager_inst.add_one_monitor(fifo_monitor_2313);
    sample_manager_inst.add_one_monitor(fifo_monitor_2314);
    sample_manager_inst.add_one_monitor(fifo_monitor_2315);
    sample_manager_inst.add_one_monitor(fifo_monitor_2316);
    sample_manager_inst.add_one_monitor(fifo_monitor_2317);
    sample_manager_inst.add_one_monitor(fifo_monitor_2318);
    sample_manager_inst.add_one_monitor(fifo_monitor_2319);
    sample_manager_inst.add_one_monitor(fifo_monitor_2320);
    sample_manager_inst.add_one_monitor(fifo_monitor_2321);
    sample_manager_inst.add_one_monitor(fifo_monitor_2322);
    sample_manager_inst.add_one_monitor(fifo_monitor_2323);
    sample_manager_inst.add_one_monitor(fifo_monitor_2324);
    sample_manager_inst.add_one_monitor(fifo_monitor_2325);
    sample_manager_inst.add_one_monitor(fifo_monitor_2326);
    sample_manager_inst.add_one_monitor(fifo_monitor_2327);
    sample_manager_inst.add_one_monitor(fifo_monitor_2328);
    sample_manager_inst.add_one_monitor(fifo_monitor_2329);
    sample_manager_inst.add_one_monitor(fifo_monitor_2330);
    sample_manager_inst.add_one_monitor(fifo_monitor_2331);
    sample_manager_inst.add_one_monitor(fifo_monitor_2332);
    sample_manager_inst.add_one_monitor(fifo_monitor_2333);
    sample_manager_inst.add_one_monitor(fifo_monitor_2334);
    sample_manager_inst.add_one_monitor(fifo_monitor_2335);
    sample_manager_inst.add_one_monitor(fifo_monitor_2336);
    sample_manager_inst.add_one_monitor(fifo_monitor_2337);
    sample_manager_inst.add_one_monitor(fifo_monitor_2338);
    sample_manager_inst.add_one_monitor(fifo_monitor_2339);
    sample_manager_inst.add_one_monitor(fifo_monitor_2340);
    sample_manager_inst.add_one_monitor(fifo_monitor_2341);
    sample_manager_inst.add_one_monitor(fifo_monitor_2342);
    sample_manager_inst.add_one_monitor(fifo_monitor_2343);
    sample_manager_inst.add_one_monitor(fifo_monitor_2344);
    sample_manager_inst.add_one_monitor(fifo_monitor_2345);
    sample_manager_inst.add_one_monitor(fifo_monitor_2346);
    sample_manager_inst.add_one_monitor(fifo_monitor_2347);
    sample_manager_inst.add_one_monitor(fifo_monitor_2348);
    sample_manager_inst.add_one_monitor(fifo_monitor_2349);
    sample_manager_inst.add_one_monitor(fifo_monitor_2350);
    sample_manager_inst.add_one_monitor(fifo_monitor_2351);
    sample_manager_inst.add_one_monitor(fifo_monitor_2352);
    sample_manager_inst.add_one_monitor(fifo_monitor_2353);
    sample_manager_inst.add_one_monitor(fifo_monitor_2354);
    sample_manager_inst.add_one_monitor(fifo_monitor_2355);
    sample_manager_inst.add_one_monitor(fifo_monitor_2356);
    sample_manager_inst.add_one_monitor(fifo_monitor_2357);
    sample_manager_inst.add_one_monitor(fifo_monitor_2358);
    sample_manager_inst.add_one_monitor(fifo_monitor_2359);
    sample_manager_inst.add_one_monitor(fifo_monitor_2360);
    sample_manager_inst.add_one_monitor(fifo_monitor_2361);
    sample_manager_inst.add_one_monitor(fifo_monitor_2362);
    sample_manager_inst.add_one_monitor(fifo_monitor_2363);
    sample_manager_inst.add_one_monitor(fifo_monitor_2364);
    sample_manager_inst.add_one_monitor(fifo_monitor_2365);
    sample_manager_inst.add_one_monitor(fifo_monitor_2366);
    sample_manager_inst.add_one_monitor(fifo_monitor_2367);
    sample_manager_inst.add_one_monitor(fifo_monitor_2368);
    sample_manager_inst.add_one_monitor(fifo_monitor_2369);
    sample_manager_inst.add_one_monitor(fifo_monitor_2370);
    sample_manager_inst.add_one_monitor(fifo_monitor_2371);
    sample_manager_inst.add_one_monitor(fifo_monitor_2372);
    sample_manager_inst.add_one_monitor(fifo_monitor_2373);
    sample_manager_inst.add_one_monitor(fifo_monitor_2374);
    sample_manager_inst.add_one_monitor(fifo_monitor_2375);
    sample_manager_inst.add_one_monitor(fifo_monitor_2376);
    sample_manager_inst.add_one_monitor(fifo_monitor_2377);
    sample_manager_inst.add_one_monitor(fifo_monitor_2378);
    sample_manager_inst.add_one_monitor(fifo_monitor_2379);
    sample_manager_inst.add_one_monitor(fifo_monitor_2380);
    sample_manager_inst.add_one_monitor(fifo_monitor_2381);
    sample_manager_inst.add_one_monitor(fifo_monitor_2382);
    sample_manager_inst.add_one_monitor(fifo_monitor_2383);
    sample_manager_inst.add_one_monitor(fifo_monitor_2384);
    sample_manager_inst.add_one_monitor(fifo_monitor_2385);
    sample_manager_inst.add_one_monitor(fifo_monitor_2386);
    sample_manager_inst.add_one_monitor(fifo_monitor_2387);
    sample_manager_inst.add_one_monitor(fifo_monitor_2388);
    sample_manager_inst.add_one_monitor(fifo_monitor_2389);
    sample_manager_inst.add_one_monitor(fifo_monitor_2390);
    sample_manager_inst.add_one_monitor(fifo_monitor_2391);
    sample_manager_inst.add_one_monitor(fifo_monitor_2392);
    sample_manager_inst.add_one_monitor(fifo_monitor_2393);
    sample_manager_inst.add_one_monitor(fifo_monitor_2394);
    sample_manager_inst.add_one_monitor(fifo_monitor_2395);
    sample_manager_inst.add_one_monitor(fifo_monitor_2396);
    sample_manager_inst.add_one_monitor(fifo_monitor_2397);
    sample_manager_inst.add_one_monitor(fifo_monitor_2398);
    sample_manager_inst.add_one_monitor(fifo_monitor_2399);
    sample_manager_inst.add_one_monitor(fifo_monitor_2400);
    sample_manager_inst.add_one_monitor(fifo_monitor_2401);
    sample_manager_inst.add_one_monitor(fifo_monitor_2402);
    sample_manager_inst.add_one_monitor(fifo_monitor_2403);
    sample_manager_inst.add_one_monitor(fifo_monitor_2404);
    sample_manager_inst.add_one_monitor(fifo_monitor_2405);
    sample_manager_inst.add_one_monitor(fifo_monitor_2406);
    sample_manager_inst.add_one_monitor(fifo_monitor_2407);
    sample_manager_inst.add_one_monitor(fifo_monitor_2408);
    sample_manager_inst.add_one_monitor(fifo_monitor_2409);
    sample_manager_inst.add_one_monitor(fifo_monitor_2410);
    sample_manager_inst.add_one_monitor(fifo_monitor_2411);
    sample_manager_inst.add_one_monitor(fifo_monitor_2412);
    sample_manager_inst.add_one_monitor(fifo_monitor_2413);
    sample_manager_inst.add_one_monitor(fifo_monitor_2414);
    sample_manager_inst.add_one_monitor(fifo_monitor_2415);
    sample_manager_inst.add_one_monitor(fifo_monitor_2416);
    sample_manager_inst.add_one_monitor(fifo_monitor_2417);
    sample_manager_inst.add_one_monitor(fifo_monitor_2418);
    sample_manager_inst.add_one_monitor(fifo_monitor_2419);
    sample_manager_inst.add_one_monitor(fifo_monitor_2420);
    sample_manager_inst.add_one_monitor(fifo_monitor_2421);
    sample_manager_inst.add_one_monitor(fifo_monitor_2422);
    sample_manager_inst.add_one_monitor(fifo_monitor_2423);
    sample_manager_inst.add_one_monitor(fifo_monitor_2424);
    sample_manager_inst.add_one_monitor(fifo_monitor_2425);
    sample_manager_inst.add_one_monitor(fifo_monitor_2426);
    sample_manager_inst.add_one_monitor(fifo_monitor_2427);
    sample_manager_inst.add_one_monitor(fifo_monitor_2428);
    sample_manager_inst.add_one_monitor(fifo_monitor_2429);
    sample_manager_inst.add_one_monitor(fifo_monitor_2430);
    sample_manager_inst.add_one_monitor(fifo_monitor_2431);
    sample_manager_inst.add_one_monitor(fifo_monitor_2432);
    sample_manager_inst.add_one_monitor(fifo_monitor_2433);
    sample_manager_inst.add_one_monitor(fifo_monitor_2434);
    sample_manager_inst.add_one_monitor(fifo_monitor_2435);
    sample_manager_inst.add_one_monitor(fifo_monitor_2436);
    sample_manager_inst.add_one_monitor(fifo_monitor_2437);
    sample_manager_inst.add_one_monitor(fifo_monitor_2438);
    sample_manager_inst.add_one_monitor(fifo_monitor_2439);
    sample_manager_inst.add_one_monitor(fifo_monitor_2440);
    sample_manager_inst.add_one_monitor(fifo_monitor_2441);
    sample_manager_inst.add_one_monitor(fifo_monitor_2442);
    sample_manager_inst.add_one_monitor(fifo_monitor_2443);
    sample_manager_inst.add_one_monitor(fifo_monitor_2444);
    sample_manager_inst.add_one_monitor(fifo_monitor_2445);
    sample_manager_inst.add_one_monitor(fifo_monitor_2446);
    sample_manager_inst.add_one_monitor(fifo_monitor_2447);
    sample_manager_inst.add_one_monitor(fifo_monitor_2448);
    sample_manager_inst.add_one_monitor(fifo_monitor_2449);
    sample_manager_inst.add_one_monitor(fifo_monitor_2450);
    sample_manager_inst.add_one_monitor(fifo_monitor_2451);
    sample_manager_inst.add_one_monitor(fifo_monitor_2452);
    sample_manager_inst.add_one_monitor(fifo_monitor_2453);
    sample_manager_inst.add_one_monitor(fifo_monitor_2454);
    sample_manager_inst.add_one_monitor(fifo_monitor_2455);
    sample_manager_inst.add_one_monitor(fifo_monitor_2456);
    sample_manager_inst.add_one_monitor(fifo_monitor_2457);
    sample_manager_inst.add_one_monitor(fifo_monitor_2458);
    sample_manager_inst.add_one_monitor(fifo_monitor_2459);
    sample_manager_inst.add_one_monitor(fifo_monitor_2460);
    sample_manager_inst.add_one_monitor(fifo_monitor_2461);
    sample_manager_inst.add_one_monitor(fifo_monitor_2462);
    sample_manager_inst.add_one_monitor(fifo_monitor_2463);
    sample_manager_inst.add_one_monitor(fifo_monitor_2464);
    sample_manager_inst.add_one_monitor(fifo_monitor_2465);
    sample_manager_inst.add_one_monitor(fifo_monitor_2466);
    sample_manager_inst.add_one_monitor(fifo_monitor_2467);
    sample_manager_inst.add_one_monitor(fifo_monitor_2468);
    sample_manager_inst.add_one_monitor(fifo_monitor_2469);
    sample_manager_inst.add_one_monitor(fifo_monitor_2470);
    sample_manager_inst.add_one_monitor(fifo_monitor_2471);
    sample_manager_inst.add_one_monitor(fifo_monitor_2472);
    sample_manager_inst.add_one_monitor(fifo_monitor_2473);
    sample_manager_inst.add_one_monitor(fifo_monitor_2474);
    sample_manager_inst.add_one_monitor(fifo_monitor_2475);
    sample_manager_inst.add_one_monitor(fifo_monitor_2476);
    sample_manager_inst.add_one_monitor(fifo_monitor_2477);
    sample_manager_inst.add_one_monitor(fifo_monitor_2478);
    sample_manager_inst.add_one_monitor(fifo_monitor_2479);
    sample_manager_inst.add_one_monitor(fifo_monitor_2480);
    sample_manager_inst.add_one_monitor(fifo_monitor_2481);
    sample_manager_inst.add_one_monitor(fifo_monitor_2482);
    sample_manager_inst.add_one_monitor(fifo_monitor_2483);
    sample_manager_inst.add_one_monitor(fifo_monitor_2484);
    sample_manager_inst.add_one_monitor(fifo_monitor_2485);
    sample_manager_inst.add_one_monitor(fifo_monitor_2486);
    sample_manager_inst.add_one_monitor(fifo_monitor_2487);
    sample_manager_inst.add_one_monitor(fifo_monitor_2488);
    sample_manager_inst.add_one_monitor(fifo_monitor_2489);
    sample_manager_inst.add_one_monitor(fifo_monitor_2490);
    sample_manager_inst.add_one_monitor(fifo_monitor_2491);
    sample_manager_inst.add_one_monitor(fifo_monitor_2492);
    sample_manager_inst.add_one_monitor(fifo_monitor_2493);
    sample_manager_inst.add_one_monitor(fifo_monitor_2494);
    sample_manager_inst.add_one_monitor(fifo_monitor_2495);
    sample_manager_inst.add_one_monitor(fifo_monitor_2496);
    sample_manager_inst.add_one_monitor(fifo_monitor_2497);
    sample_manager_inst.add_one_monitor(fifo_monitor_2498);
    sample_manager_inst.add_one_monitor(fifo_monitor_2499);
    sample_manager_inst.add_one_monitor(fifo_monitor_2500);
    sample_manager_inst.add_one_monitor(fifo_monitor_2501);
    sample_manager_inst.add_one_monitor(fifo_monitor_2502);
    sample_manager_inst.add_one_monitor(fifo_monitor_2503);
    sample_manager_inst.add_one_monitor(fifo_monitor_2504);
    sample_manager_inst.add_one_monitor(fifo_monitor_2505);
    sample_manager_inst.add_one_monitor(fifo_monitor_2506);
    sample_manager_inst.add_one_monitor(fifo_monitor_2507);
    sample_manager_inst.add_one_monitor(fifo_monitor_2508);
    sample_manager_inst.add_one_monitor(fifo_monitor_2509);
    sample_manager_inst.add_one_monitor(fifo_monitor_2510);
    sample_manager_inst.add_one_monitor(fifo_monitor_2511);
    sample_manager_inst.add_one_monitor(fifo_monitor_2512);
    sample_manager_inst.add_one_monitor(fifo_monitor_2513);
    sample_manager_inst.add_one_monitor(fifo_monitor_2514);
    sample_manager_inst.add_one_monitor(fifo_monitor_2515);
    sample_manager_inst.add_one_monitor(fifo_monitor_2516);
    sample_manager_inst.add_one_monitor(fifo_monitor_2517);
    sample_manager_inst.add_one_monitor(fifo_monitor_2518);
    sample_manager_inst.add_one_monitor(fifo_monitor_2519);
    sample_manager_inst.add_one_monitor(fifo_monitor_2520);
    sample_manager_inst.add_one_monitor(fifo_monitor_2521);
    sample_manager_inst.add_one_monitor(fifo_monitor_2522);
    sample_manager_inst.add_one_monitor(fifo_monitor_2523);
    sample_manager_inst.add_one_monitor(fifo_monitor_2524);
    sample_manager_inst.add_one_monitor(fifo_monitor_2525);
    sample_manager_inst.add_one_monitor(fifo_monitor_2526);
    sample_manager_inst.add_one_monitor(fifo_monitor_2527);
    sample_manager_inst.add_one_monitor(fifo_monitor_2528);
    sample_manager_inst.add_one_monitor(fifo_monitor_2529);
    sample_manager_inst.add_one_monitor(fifo_monitor_2530);
    sample_manager_inst.add_one_monitor(fifo_monitor_2531);
    sample_manager_inst.add_one_monitor(fifo_monitor_2532);
    sample_manager_inst.add_one_monitor(fifo_monitor_2533);
    sample_manager_inst.add_one_monitor(fifo_monitor_2534);
    sample_manager_inst.add_one_monitor(fifo_monitor_2535);
    sample_manager_inst.add_one_monitor(fifo_monitor_2536);
    sample_manager_inst.add_one_monitor(fifo_monitor_2537);
    sample_manager_inst.add_one_monitor(fifo_monitor_2538);
    sample_manager_inst.add_one_monitor(fifo_monitor_2539);
    sample_manager_inst.add_one_monitor(fifo_monitor_2540);
    sample_manager_inst.add_one_monitor(fifo_monitor_2541);
    sample_manager_inst.add_one_monitor(fifo_monitor_2542);
    sample_manager_inst.add_one_monitor(fifo_monitor_2543);
    sample_manager_inst.add_one_monitor(fifo_monitor_2544);
    sample_manager_inst.add_one_monitor(fifo_monitor_2545);
    sample_manager_inst.add_one_monitor(fifo_monitor_2546);
    sample_manager_inst.add_one_monitor(fifo_monitor_2547);
    sample_manager_inst.add_one_monitor(fifo_monitor_2548);
    sample_manager_inst.add_one_monitor(fifo_monitor_2549);
    sample_manager_inst.add_one_monitor(fifo_monitor_2550);
    sample_manager_inst.add_one_monitor(fifo_monitor_2551);
    sample_manager_inst.add_one_monitor(fifo_monitor_2552);
    sample_manager_inst.add_one_monitor(fifo_monitor_2553);
    sample_manager_inst.add_one_monitor(fifo_monitor_2554);
    sample_manager_inst.add_one_monitor(fifo_monitor_2555);
    sample_manager_inst.add_one_monitor(fifo_monitor_2556);
    sample_manager_inst.add_one_monitor(fifo_monitor_2557);
    sample_manager_inst.add_one_monitor(fifo_monitor_2558);
    sample_manager_inst.add_one_monitor(fifo_monitor_2559);
    sample_manager_inst.add_one_monitor(fifo_monitor_2560);
    sample_manager_inst.add_one_monitor(fifo_monitor_2561);
    sample_manager_inst.add_one_monitor(fifo_monitor_2562);
    sample_manager_inst.add_one_monitor(fifo_monitor_2563);
    sample_manager_inst.add_one_monitor(fifo_monitor_2564);
    sample_manager_inst.add_one_monitor(fifo_monitor_2565);
    sample_manager_inst.add_one_monitor(fifo_monitor_2566);
    sample_manager_inst.add_one_monitor(fifo_monitor_2567);
    sample_manager_inst.add_one_monitor(fifo_monitor_2568);
    sample_manager_inst.add_one_monitor(fifo_monitor_2569);
    sample_manager_inst.add_one_monitor(fifo_monitor_2570);
    sample_manager_inst.add_one_monitor(fifo_monitor_2571);
    sample_manager_inst.add_one_monitor(fifo_monitor_2572);
    sample_manager_inst.add_one_monitor(fifo_monitor_2573);
    sample_manager_inst.add_one_monitor(fifo_monitor_2574);
    sample_manager_inst.add_one_monitor(fifo_monitor_2575);
    sample_manager_inst.add_one_monitor(fifo_monitor_2576);
    sample_manager_inst.add_one_monitor(fifo_monitor_2577);
    sample_manager_inst.add_one_monitor(fifo_monitor_2578);
    sample_manager_inst.add_one_monitor(fifo_monitor_2579);
    sample_manager_inst.add_one_monitor(fifo_monitor_2580);
    sample_manager_inst.add_one_monitor(fifo_monitor_2581);
    sample_manager_inst.add_one_monitor(fifo_monitor_2582);
    sample_manager_inst.add_one_monitor(fifo_monitor_2583);
    sample_manager_inst.add_one_monitor(fifo_monitor_2584);
    sample_manager_inst.add_one_monitor(fifo_monitor_2585);
    sample_manager_inst.add_one_monitor(fifo_monitor_2586);
    sample_manager_inst.add_one_monitor(fifo_monitor_2587);
    sample_manager_inst.add_one_monitor(fifo_monitor_2588);
    sample_manager_inst.add_one_monitor(fifo_monitor_2589);
    sample_manager_inst.add_one_monitor(fifo_monitor_2590);
    sample_manager_inst.add_one_monitor(fifo_monitor_2591);
    sample_manager_inst.add_one_monitor(fifo_monitor_2592);
    sample_manager_inst.add_one_monitor(fifo_monitor_2593);
    sample_manager_inst.add_one_monitor(fifo_monitor_2594);
    sample_manager_inst.add_one_monitor(fifo_monitor_2595);
    sample_manager_inst.add_one_monitor(fifo_monitor_2596);
    sample_manager_inst.add_one_monitor(fifo_monitor_2597);
    sample_manager_inst.add_one_monitor(fifo_monitor_2598);
    sample_manager_inst.add_one_monitor(fifo_monitor_2599);
    sample_manager_inst.add_one_monitor(fifo_monitor_2600);
    sample_manager_inst.add_one_monitor(fifo_monitor_2601);
    sample_manager_inst.add_one_monitor(fifo_monitor_2602);
    sample_manager_inst.add_one_monitor(fifo_monitor_2603);
    sample_manager_inst.add_one_monitor(fifo_monitor_2604);
    sample_manager_inst.add_one_monitor(fifo_monitor_2605);
    sample_manager_inst.add_one_monitor(fifo_monitor_2606);
    sample_manager_inst.add_one_monitor(fifo_monitor_2607);
    sample_manager_inst.add_one_monitor(fifo_monitor_2608);
    sample_manager_inst.add_one_monitor(fifo_monitor_2609);
    sample_manager_inst.add_one_monitor(fifo_monitor_2610);
    sample_manager_inst.add_one_monitor(fifo_monitor_2611);
    sample_manager_inst.add_one_monitor(fifo_monitor_2612);
    sample_manager_inst.add_one_monitor(fifo_monitor_2613);
    sample_manager_inst.add_one_monitor(fifo_monitor_2614);
    sample_manager_inst.add_one_monitor(fifo_monitor_2615);
    sample_manager_inst.add_one_monitor(fifo_monitor_2616);
    sample_manager_inst.add_one_monitor(fifo_monitor_2617);
    sample_manager_inst.add_one_monitor(fifo_monitor_2618);
    sample_manager_inst.add_one_monitor(fifo_monitor_2619);
    sample_manager_inst.add_one_monitor(fifo_monitor_2620);
    sample_manager_inst.add_one_monitor(fifo_monitor_2621);
    sample_manager_inst.add_one_monitor(fifo_monitor_2622);
    sample_manager_inst.add_one_monitor(fifo_monitor_2623);
    sample_manager_inst.add_one_monitor(fifo_monitor_2624);
    sample_manager_inst.add_one_monitor(fifo_monitor_2625);
    sample_manager_inst.add_one_monitor(fifo_monitor_2626);
    sample_manager_inst.add_one_monitor(fifo_monitor_2627);
    sample_manager_inst.add_one_monitor(fifo_monitor_2628);
    sample_manager_inst.add_one_monitor(fifo_monitor_2629);
    sample_manager_inst.add_one_monitor(fifo_monitor_2630);
    sample_manager_inst.add_one_monitor(fifo_monitor_2631);
    sample_manager_inst.add_one_monitor(fifo_monitor_2632);
    sample_manager_inst.add_one_monitor(fifo_monitor_2633);
    sample_manager_inst.add_one_monitor(fifo_monitor_2634);
    sample_manager_inst.add_one_monitor(fifo_monitor_2635);
    sample_manager_inst.add_one_monitor(fifo_monitor_2636);
    sample_manager_inst.add_one_monitor(fifo_monitor_2637);
    sample_manager_inst.add_one_monitor(fifo_monitor_2638);
    sample_manager_inst.add_one_monitor(fifo_monitor_2639);
    sample_manager_inst.add_one_monitor(fifo_monitor_2640);
    sample_manager_inst.add_one_monitor(fifo_monitor_2641);
    sample_manager_inst.add_one_monitor(fifo_monitor_2642);
    sample_manager_inst.add_one_monitor(fifo_monitor_2643);
    sample_manager_inst.add_one_monitor(fifo_monitor_2644);
    sample_manager_inst.add_one_monitor(fifo_monitor_2645);
    sample_manager_inst.add_one_monitor(fifo_monitor_2646);
    sample_manager_inst.add_one_monitor(fifo_monitor_2647);
    sample_manager_inst.add_one_monitor(fifo_monitor_2648);
    sample_manager_inst.add_one_monitor(fifo_monitor_2649);
    sample_manager_inst.add_one_monitor(fifo_monitor_2650);
    sample_manager_inst.add_one_monitor(fifo_monitor_2651);
    sample_manager_inst.add_one_monitor(fifo_monitor_2652);
    sample_manager_inst.add_one_monitor(fifo_monitor_2653);
    sample_manager_inst.add_one_monitor(fifo_monitor_2654);
    sample_manager_inst.add_one_monitor(fifo_monitor_2655);
    sample_manager_inst.add_one_monitor(fifo_monitor_2656);
    sample_manager_inst.add_one_monitor(fifo_monitor_2657);
    sample_manager_inst.add_one_monitor(fifo_monitor_2658);
    sample_manager_inst.add_one_monitor(fifo_monitor_2659);
    sample_manager_inst.add_one_monitor(fifo_monitor_2660);
    sample_manager_inst.add_one_monitor(fifo_monitor_2661);
    sample_manager_inst.add_one_monitor(fifo_monitor_2662);
    sample_manager_inst.add_one_monitor(fifo_monitor_2663);
    sample_manager_inst.add_one_monitor(fifo_monitor_2664);
    sample_manager_inst.add_one_monitor(fifo_monitor_2665);
    sample_manager_inst.add_one_monitor(fifo_monitor_2666);
    sample_manager_inst.add_one_monitor(fifo_monitor_2667);
    sample_manager_inst.add_one_monitor(fifo_monitor_2668);
    sample_manager_inst.add_one_monitor(fifo_monitor_2669);
    sample_manager_inst.add_one_monitor(fifo_monitor_2670);
    sample_manager_inst.add_one_monitor(fifo_monitor_2671);
    sample_manager_inst.add_one_monitor(fifo_monitor_2672);
    sample_manager_inst.add_one_monitor(fifo_monitor_2673);
    sample_manager_inst.add_one_monitor(fifo_monitor_2674);
    sample_manager_inst.add_one_monitor(fifo_monitor_2675);
    sample_manager_inst.add_one_monitor(fifo_monitor_2676);
    sample_manager_inst.add_one_monitor(fifo_monitor_2677);
    sample_manager_inst.add_one_monitor(fifo_monitor_2678);
    sample_manager_inst.add_one_monitor(fifo_monitor_2679);
    sample_manager_inst.add_one_monitor(fifo_monitor_2680);
    sample_manager_inst.add_one_monitor(fifo_monitor_2681);
    sample_manager_inst.add_one_monitor(fifo_monitor_2682);
    sample_manager_inst.add_one_monitor(fifo_monitor_2683);
    sample_manager_inst.add_one_monitor(fifo_monitor_2684);
    sample_manager_inst.add_one_monitor(fifo_monitor_2685);
    sample_manager_inst.add_one_monitor(fifo_monitor_2686);
    sample_manager_inst.add_one_monitor(fifo_monitor_2687);
    sample_manager_inst.add_one_monitor(fifo_monitor_2688);
    sample_manager_inst.add_one_monitor(fifo_monitor_2689);
    sample_manager_inst.add_one_monitor(fifo_monitor_2690);
    sample_manager_inst.add_one_monitor(fifo_monitor_2691);
    sample_manager_inst.add_one_monitor(fifo_monitor_2692);
    sample_manager_inst.add_one_monitor(fifo_monitor_2693);
    sample_manager_inst.add_one_monitor(fifo_monitor_2694);
    sample_manager_inst.add_one_monitor(fifo_monitor_2695);
    sample_manager_inst.add_one_monitor(fifo_monitor_2696);
    sample_manager_inst.add_one_monitor(fifo_monitor_2697);
    sample_manager_inst.add_one_monitor(fifo_monitor_2698);
    sample_manager_inst.add_one_monitor(fifo_monitor_2699);
    sample_manager_inst.add_one_monitor(fifo_monitor_2700);
    sample_manager_inst.add_one_monitor(fifo_monitor_2701);
    sample_manager_inst.add_one_monitor(fifo_monitor_2702);
    sample_manager_inst.add_one_monitor(fifo_monitor_2703);
    sample_manager_inst.add_one_monitor(fifo_monitor_2704);
    sample_manager_inst.add_one_monitor(fifo_monitor_2705);
    sample_manager_inst.add_one_monitor(fifo_monitor_2706);
    sample_manager_inst.add_one_monitor(fifo_monitor_2707);
    sample_manager_inst.add_one_monitor(fifo_monitor_2708);
    sample_manager_inst.add_one_monitor(fifo_monitor_2709);
    sample_manager_inst.add_one_monitor(fifo_monitor_2710);
    sample_manager_inst.add_one_monitor(fifo_monitor_2711);
    sample_manager_inst.add_one_monitor(fifo_monitor_2712);
    sample_manager_inst.add_one_monitor(fifo_monitor_2713);
    sample_manager_inst.add_one_monitor(fifo_monitor_2714);
    sample_manager_inst.add_one_monitor(process_monitor_1);
    sample_manager_inst.add_one_monitor(process_monitor_2);
    sample_manager_inst.add_one_monitor(process_monitor_3);
    sample_manager_inst.add_one_monitor(process_monitor_4);
    sample_manager_inst.add_one_monitor(module_monitor_1);
    sample_manager_inst.add_one_monitor(module_monitor_2);
    sample_manager_inst.add_one_monitor(module_monitor_3);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_1);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_1);
    
    fork
        sample_manager_inst.start_monitor();
        last_transaction_done;
    join
    disable fork;

    sample_manager_inst.start_dump();
end

    task last_transaction_done();
        wait(reset == 0);
        while(1) begin
            if (finish == 1'b1) begin
                @(negedge clock);
                break;
            end
            else
                @(posedge clock);
        end
    endtask


endmodule
